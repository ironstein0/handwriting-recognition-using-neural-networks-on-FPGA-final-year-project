module ROM(
	input wire clk,
	input wire enable,
	input wire [11:0] address,
	output reg [15:0] data
	);

	reg [15:0] weights [4050:0x];

	initial begin
		weights[0] <= 0000000010001101;
		weights[1] <= 0000000101100100;
		weights[2] <= 1000010000101011;
		weights[3] <= 0000000101110010;
		weights[4] <= 0000110110101111;
		weights[5] <= 0000011101100101;
		weights[6] <= 0000010100111110;
		weights[7] <= 0000000000000001;
		weights[8] <= 1000000101010010;
		weights[9] <= 1000101111000011;
		weights[10] <= 0000011101111100;
		weights[11] <= 0000001001010110;
		weights[12] <= 1000010111111010;
		weights[13] <= 0000101010100001;
		weights[14] <= 0000000001010101;
		weights[15] <= 1000101011101110;
		weights[16] <= 0000010011101001;
		weights[17] <= 1000000001000010;
		weights[18] <= 0000100001100000;
		weights[19] <= 0000001010100101;
		weights[20] <= 0000001000100111;
		weights[21] <= 1000010101010011;
		weights[22] <= 1000011110101000;
		weights[23] <= 1000100011101000;
		weights[24] <= 0000101100111101;
		weights[25] <= 0000001000010000;
		weights[26] <= 1000100010000011;
		weights[27] <= 0000010011110000;
		weights[28] <= 0000100101111001;
		weights[29] <= 0000101011110001;
		weights[30] <= 1000101111110000;
		weights[31] <= 0000000011110101;
		weights[32] <= 1000001001000100;
		weights[33] <= 1000011010110110;
		weights[34] <= 1000001011000001;
		weights[35] <= 0000100001011011;
		weights[36] <= 0000010010100111;
		weights[37] <= 0000001001101010;
		weights[38] <= 0000010011100111;
		weights[39] <= 0000111001010011;
		weights[40] <= 1000101000101010;
		weights[41] <= 1001010100000001;
		weights[42] <= 0001000010001010;
		weights[43] <= 1000010011110011;
		weights[44] <= 0000101111011101;
		weights[45] <= 1000000100011010;
		weights[46] <= 1000000110010010;
		weights[47] <= 1000011001001001;
		weights[48] <= 0000110011110101;
		weights[49] <= 1000100100101110;
		weights[50] <= 0000101111011111;
		weights[51] <= 0000001000001011;
		weights[52] <= 1000000010001011;
		weights[53] <= 0000100010001101;
		weights[54] <= 1000101001100001;
		weights[55] <= 0001000000011110;
		weights[56] <= 1000000010011101;
		weights[57] <= 0000111110011000;
		weights[58] <= 1000010111011000;
		weights[59] <= 0000010011011101;
		weights[60] <= 1000001110011100;
		weights[61] <= 0000001000011101;
		weights[62] <= 0000100001110011;
		weights[63] <= 1000010001000001;
		weights[64] <= 1001000001000000;
		weights[65] <= 1001001011011100;
		weights[66] <= 1000000011010110;
		weights[67] <= 1000001010011001;
		weights[68] <= 1001011110100010;
		weights[69] <= 1000110110111101;
		weights[70] <= 1000100000001100;
		weights[71] <= 1000001100010010;
		weights[72] <= 0000100110001100;
		weights[73] <= 1000011010010101;
		weights[74] <= 1000000000111110;
		weights[75] <= 1000011010100011;
		weights[76] <= 1000000000010101;
		weights[77] <= 1000011111110000;
		weights[78] <= 1000010010100101;
		weights[79] <= 1000000000000001;
		weights[80] <= 1000011101111000;
		weights[81] <= 1000001110111101;
		weights[82] <= 0000001111001111;
		weights[83] <= 1000010011011001;
		weights[84] <= 1000001111001101;
		weights[85] <= 1000010101000000;
		weights[86] <= 1000110111001101;
		weights[87] <= 1000100000101001;
		weights[88] <= 0000011001111000;
		weights[89] <= 0000010010101011;
		weights[90] <= 1000001100110110;
		weights[91] <= 0000000100000001;
		weights[92] <= 1000010110000010;
		weights[93] <= 0000001110110001;
		weights[94] <= 1000000001111110;
		weights[95] <= 1000110001010110;
		weights[96] <= 1000011010111110;
		weights[97] <= 1000010111111101;
		weights[98] <= 1000011000111100;
		weights[99] <= 1000100101100010;
		weights[100] <= 0000001000110011;
		weights[101] <= 1000100101011100;
		weights[102] <= 0000000011111100;
		weights[103] <= 0000010100000000;
		weights[104] <= 0000001011111001;
		weights[105] <= 0000000100010111;
		weights[106] <= 0000000110000100;
		weights[107] <= 1000100011000101;
		weights[108] <= 0000000010010101;
		weights[109] <= 1000011001110011;
		weights[110] <= 0000000001110101;
		weights[111] <= 0001001010101001;
		weights[112] <= 0000001011010001;
		weights[113] <= 1000111101110010;
		weights[114] <= 0000000011011000;
		weights[115] <= 1000101000100110;
		weights[116] <= 1001001001110101;
		weights[117] <= 0000000100010010;
		weights[118] <= 0000000001000110;
		weights[119] <= 1000111100101110;
		weights[120] <= 1000011010101000;
		weights[121] <= 0000011100111110;
		weights[122] <= 1000011000001001;
		weights[123] <= 0000100010011011;
		weights[124] <= 0000100100011100;
		weights[125] <= 0000000001010010;
		weights[126] <= 0000110100000010;
		weights[127] <= 0000001001011101;
		weights[128] <= 0000100111100111;
		weights[129] <= 0000001110111000;
		weights[130] <= 0000010001100101;
		weights[131] <= 1000110001011110;
		weights[132] <= 0000000010101101;
		weights[133] <= 1000001010100011;
		weights[134] <= 0000001110010000;
		weights[135] <= 0000011011111110;
		weights[136] <= 0000000001100100;
		weights[137] <= 1000010010001100;
		weights[138] <= 1000001101110001;
		weights[139] <= 1000000101000100;
		weights[140] <= 1000111001101011;
		weights[141] <= 1000011110000001;
		weights[142] <= 0000100100111001;
		weights[143] <= 1000100101111000;
		weights[144] <= 1000100001101110;
		weights[145] <= 1000110001001110;
		weights[146] <= 0000101000011011;
		weights[147] <= 0000001010110011;
		weights[148] <= 1000110100100000;
		weights[149] <= 0000110110010000;
		weights[150] <= 1000010001011111;
		weights[151] <= 0000110001110111;
		weights[152] <= 1000011100011100;
		weights[153] <= 0000000010101100;
		weights[154] <= 1000000000111010;
		weights[155] <= 1000000011101100;
		weights[156] <= 0000011100110001;
		weights[157] <= 0000011001001111;
		weights[158] <= 1000010101000011;
		weights[159] <= 1000001100011101;
		weights[160] <= 0000010101010101;
		weights[161] <= 1000001100110110;
		weights[162] <= 1000000110010111;
		weights[163] <= 0000000010011011;
		weights[164] <= 1000010010110101;
		weights[165] <= 1000011110110010;
		weights[166] <= 0000100010101100;
		weights[167] <= 0000000100101000;
		weights[168] <= 0000101100000111;
		weights[169] <= 0000110000111011;
		weights[170] <= 1000011001111000;
		weights[171] <= 0000000111111110;
		weights[172] <= 0000001010011110;
		weights[173] <= 1000110100111010;
		weights[174] <= 0000000111110010;
		weights[175] <= 0000101000000100;
		weights[176] <= 1000010000101101;
		weights[177] <= 0000100100010011;
		weights[178] <= 0000011110100100;
		weights[179] <= 0000001000001010;
		weights[180] <= 0000011111011010;
		weights[181] <= 1000011001010100;
		weights[182] <= 1000111110000100;
		weights[183] <= 1000010000110110;
		weights[184] <= 0000010000000111;
		weights[185] <= 0000010100100001;
		weights[186] <= 0000001101100010;
		weights[187] <= 0000001000011000;
		weights[188] <= 0000111000001110;
		weights[189] <= 1000001111001001;
		weights[190] <= 0000001110010100;
		weights[191] <= 0000110101011001;
		weights[192] <= 1000010100000001;
		weights[193] <= 0000011010011111;
		weights[194] <= 0000011101110111;
		weights[195] <= 0000001000111111;
		weights[196] <= 0000000100000011;
		weights[197] <= 1001000100000101;
		weights[198] <= 1001001100100001;
		weights[199] <= 0000011000100011;
		weights[200] <= 1001001100100011;
		weights[201] <= 0000001101011011;
		weights[202] <= 1000000110111000;
		weights[203] <= 0000010110111111;
		weights[204] <= 1000000000010000;
		weights[205] <= 1000010010001101;
		weights[206] <= 0000110011100000;
		weights[207] <= 1000001000010101;
		weights[208] <= 0000001011110011;
		weights[209] <= 1000110001000110;
		weights[210] <= 1000011111010000;
		weights[211] <= 0000010101011000;
		weights[212] <= 0001001111100001;
		weights[213] <= 1000000111110100;
		weights[214] <= 1000011011011010;
		weights[215] <= 0000100001110001;
		weights[216] <= 1000011010100110;
		weights[217] <= 0000110100000000;
		weights[218] <= 0000101111011011;
		weights[219] <= 0000010000001000;
		weights[220] <= 0000110010001011;
		weights[221] <= 1000101110010010;
		weights[222] <= 1000101110111111;
		weights[223] <= 0000011011000110;
		weights[224] <= 1000000110010000;
		weights[225] <= 1000001101110100;
		weights[226] <= 0000001010101111;
		weights[227] <= 0000010111011100;
		weights[228] <= 0000100001000100;
		weights[229] <= 0000011101011101;
		weights[230] <= 0000101001110110;
		weights[231] <= 0000000101011101;
		weights[232] <= 0000011011000001;
		weights[233] <= 0000010101010011;
		weights[234] <= 1000100000001111;
		weights[235] <= 0000101101001011;
		weights[236] <= 1000010100011111;
		weights[237] <= 1000010010010001;
		weights[238] <= 0000110010011100;
		weights[239] <= 0000110001111000;
		weights[240] <= 1001000110101111;
		weights[241] <= 0000100101010110;
		weights[242] <= 0000101011010010;
		weights[243] <= 0000101110100101;
		weights[244] <= 1000101000101111;
		weights[245] <= 0000010001100010;
		weights[246] <= 1000000110011001;
		weights[247] <= 0000101010100110;
		weights[248] <= 1000000110001100;
		weights[249] <= 0000101110000001;
		weights[250] <= 0000100010100111;
		weights[251] <= 0000001000100011;
		weights[252] <= 0000010010000000;
		weights[253] <= 0000001011111001;
		weights[254] <= 1000110101101011;
		weights[255] <= 1000001111101000;
		weights[256] <= 1000100111100110;
		weights[257] <= 0000010010101010;
		weights[258] <= 0000000110000000;
		weights[259] <= 1000010111000011;
		weights[260] <= 0000011110100010;
		weights[261] <= 0000011111000001;
		weights[262] <= 1000010001001110;
		weights[263] <= 1000000001001100;
		weights[264] <= 0000001001101110;
		weights[265] <= 0000010011101000;
		weights[266] <= 0000011100010000;
		weights[267] <= 1000001101011000;
		weights[268] <= 0000100011100111;
		weights[269] <= 1000000100000011;
		weights[270] <= 0000101100110110;
		weights[271] <= 0000010000101110;
		weights[272] <= 1000001000000101;
		weights[273] <= 1000110000101000;
		weights[274] <= 0000001010100011;
		weights[275] <= 0000000011100110;
		weights[276] <= 0000010001110111;
		weights[277] <= 1000000010110101;
		weights[278] <= 0000000011000111;
		weights[279] <= 1000001001010001;
		weights[280] <= 0000010110100110;
		weights[281] <= 0000010001011110;
		weights[282] <= 0000111111110010;
		weights[283] <= 0000110001110001;
		weights[284] <= 1000010110111010;
		weights[285] <= 1000011010101011;
		weights[286] <= 0000010001111011;
		weights[287] <= 1000001011100000;
		weights[288] <= 1000010011101100;
		weights[289] <= 1000001101001000;
		weights[290] <= 0000100110000011;
		weights[291] <= 0000110000001011;
		weights[292] <= 1000001010111001;
		weights[293] <= 0001000001110111;
		weights[294] <= 0000110010101010;
		weights[295] <= 1000010101110110;
		weights[296] <= 1000101111101111;
		weights[297] <= 1000010110001001;
		weights[298] <= 1000100101010001;
		weights[299] <= 0000011100100000;
		weights[300] <= 1000001000111001;
		weights[301] <= 1000110010100011;
		weights[302] <= 1000100001011111;
		weights[303] <= 1001001110111111;
		weights[304] <= 1000011001010101;
		weights[305] <= 1000101110011000;
		weights[306] <= 1000100100010100;
		weights[307] <= 1000010100101101;
		weights[308] <= 1000010100111011;
		weights[309] <= 1000101011100110;
		weights[310] <= 0000010101101010;
		weights[311] <= 1000000011001000;
		weights[312] <= 0000111100101001;
		weights[313] <= 0000010111000011;
		weights[314] <= 1000101011001111;
		weights[315] <= 0000000001001010;
		weights[316] <= 0000011000010100;
		weights[317] <= 0000001000110011;
		weights[318] <= 0000110110110101;
		weights[319] <= 0000000101010000;
		weights[320] <= 0000011100100011;
		weights[321] <= 1000000110001001;
		weights[322] <= 0000010110111010;
		weights[323] <= 1000000100010110;
		weights[324] <= 1000000101010000;
		weights[325] <= 0000000110011011;
		weights[326] <= 0000001000000001;
		weights[327] <= 0000101101101111;
		weights[328] <= 0000100100101111;
		weights[329] <= 0000101000011011;
		weights[330] <= 0000001101010101;
		weights[331] <= 1000101001001010;
		weights[332] <= 1000000101000010;
		weights[333] <= 1000010110100101;
		weights[334] <= 1000110100111111;
		weights[335] <= 0000100010100010;
		weights[336] <= 0000001101110001;
		weights[337] <= 1000110111110001;
		weights[338] <= 1000110001111110;
		weights[339] <= 0000000100001000;
		weights[340] <= 0000110101000011;
		weights[341] <= 1000000001101011;
		weights[342] <= 0000010000010010;
		weights[343] <= 0000100010110011;
		weights[344] <= 0000000110000010;
		weights[345] <= 1000001101011111;
		weights[346] <= 1000110000111011;
		weights[347] <= 1000111000111010;
		weights[348] <= 0000000110001001;
		weights[349] <= 1000111000110110;
		weights[350] <= 0000000010000111;
		weights[351] <= 1000010110001011;
		weights[352] <= 1000000010100100;
		weights[353] <= 0000001011010001;
		weights[354] <= 0000001000010011;
		weights[355] <= 1000101010001111;
		weights[356] <= 1000010000000111;
		weights[357] <= 1000100000011100;
		weights[358] <= 1000011011111000;
		weights[359] <= 0000100100001001;
		weights[360] <= 1000101100001011;
		weights[361] <= 0000100010111000;
		weights[362] <= 0000000101000000;
		weights[363] <= 1000011110011010;
		weights[364] <= 1000100010010100;
		weights[365] <= 1001000001001010;
		weights[366] <= 0000101111001010;
		weights[367] <= 1001000010100111;
		weights[368] <= 1000101000000000;
		weights[369] <= 1000000100011100;
		weights[370] <= 1000001001000011;
		weights[371] <= 1000011001100000;
		weights[372] <= 1000011010001111;
		weights[373] <= 0000101010100111;
		weights[374] <= 1000001110011000;
		weights[375] <= 0000001100110011;
		weights[376] <= 1000000011110001;
		weights[377] <= 0000111101101011;
		weights[378] <= 1000110001111011;
		weights[379] <= 0000010011111011;
		weights[380] <= 0000001101100000;
		weights[381] <= 0000000011111100;
		weights[382] <= 1001000011110010;
		weights[383] <= 1000000001101110;
		weights[384] <= 1000001110000111;
		weights[385] <= 1000101111011100;
		weights[386] <= 0000100000110101;
		weights[387] <= 0000101011110110;
		weights[388] <= 0000010011000011;
		weights[389] <= 1000000010100100;
		weights[390] <= 0000000100000101;
		weights[391] <= 1000010110011010;
		weights[392] <= 1000011101001010;
		weights[393] <= 1000000011101000;
		weights[394] <= 1000011101001011;
		weights[395] <= 0000111011101011;
		weights[396] <= 1000101101011110;
		weights[397] <= 0000010110011101;
		weights[398] <= 0000010110001100;
		weights[399] <= 1000011101101101;
		weights[400] <= 0000110100101101;
		weights[401] <= 0000011101010001;
		weights[402] <= 1000000101010000;
		weights[403] <= 1000010100110010;
		weights[404] <= 0000001001110101;
		weights[405] <= 1001001111111000;
		weights[406] <= 0000110011111010;
		weights[407] <= 1000000000010000;
		weights[408] <= 1000110101000100;
		weights[409] <= 1000101100000000;
		weights[410] <= 0000010011111110;
		weights[411] <= 0000011101011100;
		weights[412] <= 0000100110110110;
		weights[413] <= 1000001110011000;
		weights[414] <= 1000000110110111;
		weights[415] <= 1000001110111111;
		weights[416] <= 1000010000010110;
		weights[417] <= 1000100110011101;
		weights[418] <= 1000000011001111;
		weights[419] <= 1000000110000011;
		weights[420] <= 1000110100001011;
		weights[421] <= 0001000100101101;
		weights[422] <= 0000010001111000;
		weights[423] <= 0000001000110111;
		weights[424] <= 0000001110111111;
		weights[425] <= 0000101100100001;
		weights[426] <= 1000000001101011;
		weights[427] <= 1001000000101111;
		weights[428] <= 0000010010101000;
		weights[429] <= 1000011111001000;
		weights[430] <= 0000010011101100;
		weights[431] <= 0000100111000110;
		weights[432] <= 0000011001101001;
		weights[433] <= 0001000101100010;
		weights[434] <= 0000000011111101;
		weights[435] <= 0000000000010110;
		weights[436] <= 1000001000111100;
		weights[437] <= 1000011010110001;
		weights[438] <= 1000010111100011;
		weights[439] <= 1000010000110001;
		weights[440] <= 1000001110011010;
		weights[441] <= 0000101100110111;
		weights[442] <= 1000101100110010;
		weights[443] <= 0000011100111010;
		weights[444] <= 0000101111100000;
		weights[445] <= 1000101000100000;
		weights[446] <= 0000000110110110;
		weights[447] <= 0000100110001011;
		weights[448] <= 1000111101110001;
		weights[449] <= 1000010000001001;
		weights[450] <= 1000110000101000;
		weights[451] <= 1001000101000100;
		weights[452] <= 0000101010011001;
		weights[453] <= 1000010010111100;
		weights[454] <= 0000100011010110;
		weights[455] <= 1000000010110011;
		weights[456] <= 1000010100010100;
		weights[457] <= 1000110000111010;
		weights[458] <= 0000110110101100;
		weights[459] <= 1000000101000010;
		weights[460] <= 0000011000011110;
		weights[461] <= 0000000001111111;
		weights[462] <= 1000000101000111;
		weights[463] <= 0000000011100110;
		weights[464] <= 1000010110010110;
		weights[465] <= 1000010010111000;
		weights[466] <= 0001010001111001;
		weights[467] <= 0000001010111010;
		weights[468] <= 1000100000011010;
		weights[469] <= 0000100001001101;
		weights[470] <= 0000000000100001;
		weights[471] <= 0000010010110001;
		weights[472] <= 1000001001100100;
		weights[473] <= 0001001101000010;
		weights[474] <= 0000010001011100;
		weights[475] <= 1000001111001001;
		weights[476] <= 1000001001101100;
		weights[477] <= 1000000011000001;
		weights[478] <= 1000000111101001;
		weights[479] <= 0000010110100101;
		weights[480] <= 0000000001110111;
		weights[481] <= 0000010001000101;
		weights[482] <= 1000100000111010;
		weights[483] <= 1000011000100111;
		weights[484] <= 1000100110011111;
		weights[485] <= 1000010101000011;
		weights[486] <= 1000101011001101;
		weights[487] <= 0000011001001111;
		weights[488] <= 1000011010111111;
		weights[489] <= 1000001111000111;
		weights[490] <= 0000110101010000;
		weights[491] <= 1000010001001001;
		weights[492] <= 0000001001111100;
		weights[493] <= 1000000110011110;
		weights[494] <= 1000000110101100;
		weights[495] <= 1000001111000000;
		weights[496] <= 0000001101000100;
		weights[497] <= 0000010100110111;
		weights[498] <= 1000100010000111;
		weights[499] <= 1000010011001001;
		weights[500] <= 0000011100110011;
		weights[501] <= 1000011100110011;
		weights[502] <= 0000010100011010;
		weights[503] <= 1000110011001010;
		weights[504] <= 0000010101000011;
		weights[505] <= 1000101011000111;
		weights[506] <= 0000000001101111;
		weights[507] <= 1000001010010011;
		weights[508] <= 1000000000101011;
		weights[509] <= 1000010101001110;
		weights[510] <= 1000001100011110;
		weights[511] <= 0000000010111011;
		weights[512] <= 0000000110000010;
		weights[513] <= 1000001110101001;
		weights[514] <= 1000001111101111;
		weights[515] <= 0000001100000110;
		weights[516] <= 0000011111110110;
		weights[517] <= 0000010000001001;
		weights[518] <= 1000000100011101;
		weights[519] <= 1000011011111101;
		weights[520] <= 1000100011111000;
		weights[521] <= 0000011001001000;
		weights[522] <= 1000110111100111;
		weights[523] <= 0000011110000110;
		weights[524] <= 1000000001110101;
		weights[525] <= 0000100000111010;
		weights[526] <= 0000001111010000;
		weights[527] <= 0000100111000110;
		weights[528] <= 0001000110001001;
		weights[529] <= 0000100000000001;
		weights[530] <= 0000010001110111;
		weights[531] <= 0000000111011011;
		weights[532] <= 0000000010111111;
		weights[533] <= 0000010000011111;
		weights[534] <= 1000010110000110;
		weights[535] <= 1000010000111100;
		weights[536] <= 0000011111000011;
		weights[537] <= 0000010100111100;
		weights[538] <= 1000111100001010;
		weights[539] <= 0000011101010100;
		weights[540] <= 0001001100100001;
		weights[541] <= 1000000101010110;
		weights[542] <= 1000000001110010;
		weights[543] <= 1000011001001000;
		weights[544] <= 0000001000000001;
		weights[545] <= 0000100111010111;
		weights[546] <= 0001001001111101;
		weights[547] <= 0010001011010000;
		weights[548] <= 0010001101000011;
		weights[549] <= 0001010111011000;
		weights[550] <= 0000100110010001;
		weights[551] <= 0000100111101101;
		weights[552] <= 0000011110100100;
		weights[553] <= 0000011110110001;
		weights[554] <= 0000000010101111;
		weights[555] <= 1000110010010000;
		weights[556] <= 0000001000001000;
		weights[557] <= 1000010010010001;
		weights[558] <= 0000011000111001;
		weights[559] <= 0000110111001110;
		weights[560] <= 0000010100010011;
		weights[561] <= 0000001001111110;
		weights[562] <= 1000010101100001;
		weights[563] <= 1000011111110010;
		weights[564] <= 1000001001010010;
		weights[565] <= 0000010000000111;
		weights[566] <= 0001001101100001;
		weights[567] <= 0000101110010110;
		weights[568] <= 0000010100010101;
		weights[569] <= 0000101001010110;
		weights[570] <= 0000011101110110;
		weights[571] <= 1000110101010111;
		weights[572] <= 0000000011000110;
		weights[573] <= 1000001111100100;
		weights[574] <= 0000101001011001;
		weights[575] <= 0000001011111111;
		weights[576] <= 0000010000001000;
		weights[577] <= 0000011000011010;
		weights[578] <= 1000011011110111;
		weights[579] <= 0000010101000101;
		weights[580] <= 1000100010010001;
		weights[581] <= 0000100011010100;
		weights[582] <= 0000000100110100;
		weights[583] <= 1000000111011010;
		weights[584] <= 0000011011111011;
		weights[585] <= 1000001000101000;
		weights[586] <= 0000100001001101;
		weights[587] <= 0000000100100010;
		weights[588] <= 1000000101000111;
		weights[589] <= 0000000011100011;
		weights[590] <= 1000000100010001;
		weights[591] <= 1000001101010000;
		weights[592] <= 1000001101110010;
		weights[593] <= 1000010000100010;
		weights[594] <= 1000000101001101;
		weights[595] <= 1000001111011111;
		weights[596] <= 0000110011111100;
		weights[597] <= 1000100100000100;
		weights[598] <= 0000000101100000;
		weights[599] <= 0000000001000101;
		weights[600] <= 1000111010010010;
		weights[601] <= 1001000101000101;
		weights[602] <= 0000101111010000;
		weights[603] <= 1000101011001000;
		weights[604] <= 1000010011110101;
		weights[605] <= 0000100110101111;
		weights[606] <= 0000000011000000;
		weights[607] <= 1000000000100111;
		weights[608] <= 0000010011100001;
		weights[609] <= 0000011110110011;
		weights[610] <= 1000010011100110;
		weights[611] <= 1000110001111010;
		weights[612] <= 1000000101101111;
		weights[613] <= 0000001011001010;
		weights[614] <= 0000001011100110;
		weights[615] <= 0000100110000110;
		weights[616] <= 0000010101011010;
		weights[617] <= 0000011011011110;
		weights[618] <= 0000010010100000;
		weights[619] <= 0000001011011011;
		weights[620] <= 0000010100001000;
		weights[621] <= 0000000011110110;
		weights[622] <= 1000010000001001;
		weights[623] <= 1000101011101100;
		weights[624] <= 1000010000010000;
		weights[625] <= 1000001010100010;
		weights[626] <= 1000011100110001;
		weights[627] <= 0000000110101011;
		weights[628] <= 1000000101001101;
		weights[629] <= 0000010110100001;
		weights[630] <= 1000000000100010;
		weights[631] <= 1000011011111110;
		weights[632] <= 1000000010100011;
		weights[633] <= 1000000001011010;
		weights[634] <= 1000001111011001;
		weights[635] <= 1000001111110111;
		weights[636] <= 1000011000010111;
		weights[637] <= 0000000010111010;
		weights[638] <= 0000001110001101;
		weights[639] <= 1000101101101110;
		weights[640] <= 1000010101010011;
		weights[641] <= 1000010110010000;
		weights[642] <= 0000000101001010;
		weights[643] <= 1000000010101001;
		weights[644] <= 0000011110111110;
		weights[645] <= 1000001000000001;
		weights[646] <= 1000010000110011;
		weights[647] <= 1000000001000000;
		weights[648] <= 0000000000101101;
		weights[649] <= 1000000010101101;
		weights[650] <= 1000001100110100;
		weights[651] <= 1000001110010101;
		weights[652] <= 0000000110111111;
		weights[653] <= 1000100011000101;
		weights[654] <= 0000000010010110;
		weights[655] <= 0000010000111010;
		weights[656] <= 1000011000111010;
		weights[657] <= 0000110101111110;
		weights[658] <= 1000110101000100;
		weights[659] <= 1000100101101011;
		weights[660] <= 0000010010101011;
		weights[661] <= 0000011110011000;
		weights[662] <= 0000000000101110;
		weights[663] <= 0000111010101101;
		weights[664] <= 0000101111011111;
		weights[665] <= 1000000101111110;
		weights[666] <= 1000011101000010;
		weights[667] <= 1000001110111001;
		weights[668] <= 1000001000011100;
		weights[669] <= 1000000101101001;
		weights[670] <= 0000000100111100;
		weights[671] <= 0000000010000111;
		weights[672] <= 1000011001000111;
		weights[673] <= 1000101011001110;
		weights[674] <= 1000100010011100;
		weights[675] <= 1001000011101100;
		weights[676] <= 1000101101100101;
		weights[677] <= 1000101010011000;
		weights[678] <= 1000100010011000;
		weights[679] <= 0000101100011111;
		weights[680] <= 0000010011010010;
		weights[681] <= 1000001000111100;
		weights[682] <= 1000100011001011;
		weights[683] <= 0000011010011011;
		weights[684] <= 1000110000000011;
		weights[685] <= 0000000010111100;
		weights[686] <= 0000101010001100;
		weights[687] <= 1000010001101011;
		weights[688] <= 1000011000001100;
		weights[689] <= 1000001111101000;
		weights[690] <= 1000011011111101;
		weights[691] <= 1000011101000100;
		weights[692] <= 1000100000011110;
		weights[693] <= 0000001011001111;
		weights[694] <= 0000000011011011;
		weights[695] <= 1000001011011110;
		weights[696] <= 1000110011101001;
		weights[697] <= 0000100011110101;
		weights[698] <= 1000001000010011;
		weights[699] <= 0000010100100111;
		weights[700] <= 0000010111100111;
		weights[701] <= 1000001000011001;
		weights[702] <= 0001000000000010;
		weights[703] <= 0000010100101100;
		weights[704] <= 1000001111011000;
		weights[705] <= 1000101111000000;
		weights[706] <= 1000000111011101;
		weights[707] <= 1000011011110110;
		weights[708] <= 1001000010001011;
		weights[709] <= 1000010111011011;
		weights[710] <= 1000110110000101;
		weights[711] <= 1000100010101100;
		weights[712] <= 1000001010101111;
		weights[713] <= 0000100001101111;
		weights[714] <= 0000011000111110;
		weights[715] <= 0001011011001011;
		weights[716] <= 1000000011001111;
		weights[717] <= 0000001001000000;
		weights[718] <= 1000101111001110;
		weights[719] <= 0000111100100000;
		weights[720] <= 0000010010010110;
		weights[721] <= 0000000001101001;
		weights[722] <= 1000001000101001;
		weights[723] <= 0000000110010101;
		weights[724] <= 1000001100111101;
		weights[725] <= 1000110001111000;
		weights[726] <= 0000010010100001;
		weights[727] <= 0000100000001000;
		weights[728] <= 1000000101100110;
		weights[729] <= 0000000110000010;
		weights[730] <= 1000011100010100;
		weights[731] <= 1000010011100001;
		weights[732] <= 1000011101011000;
		weights[733] <= 1001000001110111;
		weights[734] <= 0000011110011100;
		weights[735] <= 1000101000101100;
		weights[736] <= 1001000110100001;
		weights[737] <= 1000111101100111;
		weights[738] <= 0000110110110000;
		weights[739] <= 0000000100101011;
		weights[740] <= 0000001011111000;
		weights[741] <= 0000101100000001;
		weights[742] <= 1001000100110110;
		weights[743] <= 1000001101110010;
		weights[744] <= 1000000100000111;
		weights[745] <= 1000011000011111;
		weights[746] <= 1000000011101000;
		weights[747] <= 0000010100010110;
		weights[748] <= 0001000001010110;
		weights[749] <= 1000000101001011;
		weights[750] <= 0000011010100101;
		weights[751] <= 0000010000111000;
		weights[752] <= 0000011111000101;
		weights[753] <= 1000011110100011;
		weights[754] <= 0000001010001110;
		weights[755] <= 1000000001011010;
		weights[756] <= 1000100010010100;
		weights[757] <= 0000000100011000;
		weights[758] <= 1000011000011101;
		weights[759] <= 0000000000101110;
		weights[760] <= 1000001000101110;
		weights[761] <= 1000010101001101;
		weights[762] <= 0000001001101001;
		weights[763] <= 1000001011000101;
		weights[764] <= 0000011110111010;
		weights[765] <= 1000110001111110;
		weights[766] <= 1000011111110000;
		weights[767] <= 0000001011010100;
		weights[768] <= 0000011110100100;
		weights[769] <= 0000101111110101;
		weights[770] <= 0000011111100110;
		weights[771] <= 0000010111100111;
		weights[772] <= 1000001001000000;
		weights[773] <= 0000011000101001;
		weights[774] <= 1000001011000100;
		weights[775] <= 1000010000000111;
		weights[776] <= 0000110100111110;
		weights[777] <= 0000100111110110;
		weights[778] <= 1000101111111001;
		weights[779] <= 1000100101101000;
		weights[780] <= 1000110000011100;
		weights[781] <= 0000011001011101;
		weights[782] <= 0000001001010011;
		weights[783] <= 0000000000110101;
		weights[784] <= 1000000000111101;
		weights[785] <= 0000000011100111;
		weights[786] <= 1000011001111001;
		weights[787] <= 1000011101000000;
		weights[788] <= 0000011110001111;
		weights[789] <= 1000010011010101;
		weights[790] <= 1000100011100110;
		weights[791] <= 1000010111001010;
		weights[792] <= 0000001100011010;
		weights[793] <= 0000000000100110;
		weights[794] <= 0000000111011111;
		weights[795] <= 1000010111101100;
		weights[796] <= 0000001111000111;
		weights[797] <= 0000010010101011;
		weights[798] <= 0000011111011111;
		weights[799] <= 0000111111110000;
		weights[800] <= 1000010011010010;
		weights[801] <= 0000000011011010;
		weights[802] <= 1000101101101100;
		weights[803] <= 0000000100100011;
		weights[804] <= 1000100100011100;
		weights[805] <= 1000011001101000;
		weights[806] <= 0000100101011111;
		weights[807] <= 0000001001101100;
		weights[808] <= 1000011001110011;
		weights[809] <= 0000001111011011;
		weights[810] <= 1000000111111010;
		weights[811] <= 0000000010001101;
		weights[812] <= 1000000111001010;
		weights[813] <= 1001001010110011;
		weights[814] <= 1001001101001001;
		weights[815] <= 0000000100110100;
		weights[816] <= 1000011100010001;
		weights[817] <= 1000000100001110;
		weights[818] <= 0000011000001001;
		weights[819] <= 1000001110111001;
		weights[820] <= 1000001000000101;
		weights[821] <= 0000011001001111;
		weights[822] <= 0000001010001011;
		weights[823] <= 1000000000110001;
		weights[824] <= 1000000110000011;
		weights[825] <= 1000011011100100;
		weights[826] <= 0000101101010000;
		weights[827] <= 1000000010011101;
		weights[828] <= 1000101111011101;
		weights[829] <= 1000100110010101;
		weights[830] <= 1000011010000111;
		weights[831] <= 1000000000011000;
		weights[832] <= 1000011111011001;
		weights[833] <= 1000101111011110;
		weights[834] <= 1000010011101001;
		weights[835] <= 0000000001001001;
		weights[836] <= 1000000001011010;
		weights[837] <= 1000010010101001;
		weights[838] <= 1000000111110010;
		weights[839] <= 0000010011010110;
		weights[840] <= 0000001100111101;
		weights[841] <= 1000000001010011;
		weights[842] <= 0000000001011001;
		weights[843] <= 0000001111100010;
		weights[844] <= 0000100100001010;
		weights[845] <= 0000001100110100;
		weights[846] <= 0000000000110000;
		weights[847] <= 0000111010111101;
		weights[848] <= 1000100010010110;
		weights[849] <= 1000001111101100;
		weights[850] <= 0001000110000000;
		weights[851] <= 0000011010101110;
		weights[852] <= 1000010011111001;
		weights[853] <= 0000000011000101;
		weights[854] <= 1000001101001110;
		weights[855] <= 0000001110100100;
		weights[856] <= 0000001101001101;
		weights[857] <= 0000001010000001;
		weights[858] <= 0000010001000011;
		weights[859] <= 1000111001111110;
		weights[860] <= 1000010010001110;
		weights[861] <= 0000000101101110;
		weights[862] <= 1000011111101100;
		weights[863] <= 1000111110101111;
		weights[864] <= 0001000001000110;
		weights[865] <= 0000000101111111;
		weights[866] <= 1000010001000000;
		weights[867] <= 1000010011001110;
		weights[868] <= 0000110111001011;
		weights[869] <= 0000001011101101;
		weights[870] <= 0000110101110101;
		weights[871] <= 0000110001110000;
		weights[872] <= 1000001000101111;
		weights[873] <= 0000011001001000;
		weights[874] <= 0000011000001000;
		weights[875] <= 0000001001010001;
		weights[876] <= 0000001101111100;
		weights[877] <= 0000101101111001;
		weights[878] <= 1000111001100011;
		weights[879] <= 1000100000010101;
		weights[880] <= 1000001011110100;
		weights[881] <= 0000101100011000;
		weights[882] <= 0000001101001110;
		weights[883] <= 0000011001101111;
		weights[884] <= 0001001111011101;
		weights[885] <= 0000000110000111;
		weights[886] <= 0000001010001100;
		weights[887] <= 1000010011010111;
		weights[888] <= 0000000110011010;
		weights[889] <= 0000001101001110;
		weights[890] <= 0000011100010101;
		weights[891] <= 0000011001111111;
		weights[892] <= 1000010101110000;
		weights[893] <= 1000011010011101;
		weights[894] <= 0000010000101100;
		weights[895] <= 0000010111001000;
		weights[896] <= 1000011101000100;
		weights[897] <= 0000101100010110;
		weights[898] <= 1000001111011110;
		weights[899] <= 1000010011001001;
		weights[900] <= 0000010000100010;
		weights[901] <= 0000000111001101;
		weights[902] <= 0000100110111101;
		weights[903] <= 1000011110010011;
		weights[904] <= 1000101011101000;
		weights[905] <= 0000001100011011;
		weights[906] <= 1000010101001101;
		weights[907] <= 0000001101100011;
		weights[908] <= 1000000111010001;
		weights[909] <= 0000001010001000;
		weights[910] <= 0000010101001111;
		weights[911] <= 0000010101001010;
		weights[912] <= 0000001001000011;
		weights[913] <= 0000000100001001;
		weights[914] <= 0000000010010100;
		weights[915] <= 1000101110000100;
		weights[916] <= 1000101110011101;
		weights[917] <= 1000001010100100;
		weights[918] <= 1000000101001110;
		weights[919] <= 1000000010111100;
		weights[920] <= 0000100011100100;
		weights[921] <= 1000101001111001;
		weights[922] <= 0000001010101100;
		weights[923] <= 1000011110100010;
		weights[924] <= 1000010010111010;
		weights[925] <= 1000001101001001;
		weights[926] <= 1000010110111101;
		weights[927] <= 0000001111000110;
		weights[928] <= 0000011011110110;
		weights[929] <= 0000011000100100;
		weights[930] <= 0000010010110101;
		weights[931] <= 0000001010110000;
		weights[932] <= 1000001011011011;
		weights[933] <= 0000000000000001;
		weights[934] <= 1000001101111000;
		weights[935] <= 1000000011001100;
		weights[936] <= 1000001110011001;
		weights[937] <= 1000001010110010;
		weights[938] <= 1000010000000100;
		weights[939] <= 1000001000100101;
		weights[940] <= 0000000010001010;
		weights[941] <= 0000010101101110;
		weights[942] <= 1000001100000011;
		weights[943] <= 0001001010111000;
		weights[944] <= 1000011010001001;
		weights[945] <= 1000000011111000;
		weights[946] <= 1000011110111001;
		weights[947] <= 0000100111010000;
		weights[948] <= 0000100010000110;
		weights[949] <= 0000100111101011;
		weights[950] <= 1000000001100110;
		weights[951] <= 1000000010111001;
		weights[952] <= 0000000011101001;
		weights[953] <= 1000000100110110;
		weights[954] <= 1000010001100011;
		weights[955] <= 1000000011111010;
		weights[956] <= 0000001111010010;
		weights[957] <= 1001001101111101;
		weights[958] <= 0000010110011111;
		weights[959] <= 0000001111101000;
		weights[960] <= 0000101101110010;
		weights[961] <= 0000011111100111;
		weights[962] <= 0000111101010011;
		weights[963] <= 1000000010111110;
		weights[964] <= 1000011010000111;
		weights[965] <= 1000011001110101;
		weights[966] <= 1000000111010011;
		weights[967] <= 1000001000111100;
		weights[968] <= 0000011000110010;
		weights[969] <= 0000011111010011;
		weights[970] <= 0001100100101100;
		weights[971] <= 0001100010101011;
		weights[972] <= 0000110010010011;
		weights[973] <= 0000010111000010;
		weights[974] <= 1000001000111101;
		weights[975] <= 1000000000101111;
		weights[976] <= 1000000001001011;
		weights[977] <= 1000010000000001;
		weights[978] <= 0000000010011001;
		weights[979] <= 0000010010011110;
		weights[980] <= 0000110001100100;
		weights[981] <= 0000010000010101;
		weights[982] <= 0000111000110110;
		weights[983] <= 0000101001110001;
		weights[984] <= 0000100001111001;
		weights[985] <= 1000001111011101;
		weights[986] <= 0000011001110110;
		weights[987] <= 1000010010000010;
		weights[988] <= 1000011000011100;
		weights[989] <= 0000010101101110;
		weights[990] <= 0000111010111111;
		weights[991] <= 0001011111100000;
		weights[992] <= 0001100101010111;
		weights[993] <= 0000011110101101;
		weights[994] <= 0000000110010000;
		weights[995] <= 0000110110101000;
		weights[996] <= 0000011110110110;
		weights[997] <= 1000011100010001;
		weights[998] <= 1000010011000000;
		weights[999] <= 1000000110000110;
		weights[1000] <= 0000101111010001;
		weights[1001] <= 1000011110000011;
		weights[1002] <= 1000000000100001;
		weights[1003] <= 1000101000100011;
		weights[1004] <= 1000011001101000;
		weights[1005] <= 1000110011010101;
		weights[1006] <= 1000001011111010;
		weights[1007] <= 1000000001011110;
		weights[1008] <= 1000100101110100;
		weights[1009] <= 1000001000011000;
		weights[1010] <= 0001001001000110;
		weights[1011] <= 0000111111101010;
		weights[1012] <= 0000111000011110;
		weights[1013] <= 0000011000111000;
		weights[1014] <= 0000101010110000;
		weights[1015] <= 1000010011101010;
		weights[1016] <= 0000010110011001;
		weights[1017] <= 0000001011010111;
		weights[1018] <= 0000001000111110;
		weights[1019] <= 1000000010111100;
		weights[1020] <= 1000011010100001;
		weights[1021] <= 1000010101001101;
		weights[1022] <= 0000000010101111;
		weights[1023] <= 1000101100010100;
		weights[1024] <= 1000110001111100;
		weights[1025] <= 0000011100011100;
		weights[1026] <= 1000101001110010;
		weights[1027] <= 1000010000101110;
		weights[1028] <= 1000000110100100;
		weights[1029] <= 1000011110100000;
		weights[1030] <= 1000001111111011;
		weights[1031] <= 0000111011111011;
		weights[1032] <= 0000110101111011;
		weights[1033] <= 1000001101000110;
		weights[1034] <= 0000001101010100;
		weights[1035] <= 1000000101010010;
		weights[1036] <= 1000001011010111;
		weights[1037] <= 1000000100111001;
		weights[1038] <= 0000001101111110;
		weights[1039] <= 1000011010010110;
		weights[1040] <= 0000000101101000;
		weights[1041] <= 0000010011110101;
		weights[1042] <= 1000011011011011;
		weights[1043] <= 0000010011100111;
		weights[1044] <= 0000000000100100;
		weights[1045] <= 0000111010001110;
		weights[1046] <= 0000000011000100;
		weights[1047] <= 0000000000101001;
		weights[1048] <= 1000000010000000;
		weights[1049] <= 1000000001100110;
		weights[1050] <= 1000010001111000;
		weights[1051] <= 1000011000011001;
		weights[1052] <= 1000100000100110;
		weights[1053] <= 1000001001110101;
		weights[1054] <= 1000000001110100;
		weights[1055] <= 1000000110011011;
		weights[1056] <= 1000001100101101;
		weights[1057] <= 1001000100000101;
		weights[1058] <= 0000011001011010;
		weights[1059] <= 0000101101001000;
		weights[1060] <= 0000010010000111;
		weights[1061] <= 1000111010000101;
		weights[1062] <= 0000010111101100;
		weights[1063] <= 0000011010010011;
		weights[1064] <= 0000001000011001;
		weights[1065] <= 0001001010111100;
		weights[1066] <= 1000101000011110;
		weights[1067] <= 1000000000010110;
		weights[1068] <= 1000011010010101;
		weights[1069] <= 0000000001110001;
		weights[1070] <= 1000011001011001;
		weights[1071] <= 1000010101110110;
		weights[1072] <= 1000011010111000;
		weights[1073] <= 1000000101001001;
		weights[1074] <= 1000001111101010;
		weights[1075] <= 1000010000111111;
		weights[1076] <= 0000001000111001;
		weights[1077] <= 1000010011100101;
		weights[1078] <= 1000011110110110;
		weights[1079] <= 1000010101000000;
		weights[1080] <= 1000101111101110;
		weights[1081] <= 0000011100001001;
		weights[1082] <= 0000001010001000;
		weights[1083] <= 1000011000100010;
		weights[1084] <= 0000100001011000;
		weights[1085] <= 0000000001010101;
		weights[1086] <= 1000001010010111;
		weights[1087] <= 0000011110100011;
		weights[1088] <= 0000000000011100;
		weights[1089] <= 0000000001100111;
		weights[1090] <= 1000000010110111;
		weights[1091] <= 1000010010010010;
		weights[1092] <= 1000011111111000;
		weights[1093] <= 0000001011011100;
		weights[1094] <= 1000011111101000;
		weights[1095] <= 1000101010001111;
		weights[1096] <= 0000100000111001;
		weights[1097] <= 1000000100111011;
		weights[1098] <= 0001010110000011;
		weights[1099] <= 1001001100011110;
		weights[1100] <= 1000011010110001;
		weights[1101] <= 0000010110001000;
		weights[1102] <= 0000001001011111;
		weights[1103] <= 1000111001001111;
		weights[1104] <= 0000101101100101;
		weights[1105] <= 0000110100011101;
		weights[1106] <= 1000110110000000;
		weights[1107] <= 1000001100001011;
		weights[1108] <= 0000000100110010;
		weights[1109] <= 0000001000010101;
		weights[1110] <= 0000011011110110;
		weights[1111] <= 1000001000101110;
		weights[1112] <= 0000100011110000;
		weights[1113] <= 0000000111101010;
		weights[1114] <= 1000101101000100;
		weights[1115] <= 0000001100000101;
		weights[1116] <= 0000000110011010;
		weights[1117] <= 0000110011010111;
		weights[1118] <= 1000010101100100;
		weights[1119] <= 1000011010001000;
		weights[1120] <= 0000010000100000;
		weights[1121] <= 0000001111111111;
		weights[1122] <= 0000101100111100;
		weights[1123] <= 1000010000101010;
		weights[1124] <= 0000010101111110;
		weights[1125] <= 0000010001011011;
		weights[1126] <= 0000001100010110;
		weights[1127] <= 0000011111101000;
		weights[1128] <= 1000110101010111;
		weights[1129] <= 0000010000010110;
		weights[1130] <= 0000001000000010;
		weights[1131] <= 0000101101101100;
		weights[1132] <= 0000011100001000;
		weights[1133] <= 0000010010100011;
		weights[1134] <= 1000011110000100;
		weights[1135] <= 0000101111010010;
		weights[1136] <= 1000010101000110;
		weights[1137] <= 1000010110001001;
		weights[1138] <= 1000000100101111;
		weights[1139] <= 0000000100001101;
		weights[1140] <= 0000000001101101;
		weights[1141] <= 1000100111011001;
		weights[1142] <= 1000011110000111;
		weights[1143] <= 1000000010011111;
		weights[1144] <= 1000001101101011;
		weights[1145] <= 0000010011000000;
		weights[1146] <= 1000001001010011;
		weights[1147] <= 0000000101010100;
		weights[1148] <= 0000101001000111;
		weights[1149] <= 0000010100101010;
		weights[1150] <= 0000001010111000;
		weights[1151] <= 0000011111001010;
		weights[1152] <= 0000100000110110;
		weights[1153] <= 0000100010101110;
		weights[1154] <= 1000000011100010;
		weights[1155] <= 0000011010100100;
		weights[1156] <= 1000011111111001;
		weights[1157] <= 1000000101110110;
		weights[1158] <= 0000010011010101;
		weights[1159] <= 0000000011011101;
		weights[1160] <= 1000001010001000;
		weights[1161] <= 1000111101100101;
		weights[1162] <= 1000000111100011;
		weights[1163] <= 0000010101010010;
		weights[1164] <= 1000111011011100;
		weights[1165] <= 1000110011001001;
		weights[1166] <= 0000000000000010;
		weights[1167] <= 0000000100010000;
		weights[1168] <= 1000101100000001;
		weights[1169] <= 0000011010110011;
		weights[1170] <= 0000100001011001;
		weights[1171] <= 0000011001111010;
		weights[1172] <= 1000010100111011;
		weights[1173] <= 0000111001100100;
		weights[1174] <= 1000000110001011;
		weights[1175] <= 1000000010101101;
		weights[1176] <= 1000001100011100;
		weights[1177] <= 1000000010010011;
		weights[1178] <= 0000000100101011;
		weights[1179] <= 1000011001110110;
		weights[1180] <= 0000100000101001;
		weights[1181] <= 0000100100100001;
		weights[1182] <= 0000100010111100;
		weights[1183] <= 1000010011011011;
		weights[1184] <= 0000010000011001;
		weights[1185] <= 0001001110011100;
		weights[1186] <= 0000100100111001;
		weights[1187] <= 0000001111010000;
		weights[1188] <= 1000111110011001;
		weights[1189] <= 1000010000101010;
		weights[1190] <= 0000110010001011;
		weights[1191] <= 0001011010000010;
		weights[1192] <= 0000001101011101;
		weights[1193] <= 0000001110111110;
		weights[1194] <= 1000001010100111;
		weights[1195] <= 0000101011001110;
		weights[1196] <= 1000010101100101;
		weights[1197] <= 1000101001001110;
		weights[1198] <= 1000000001101011;
		weights[1199] <= 1000000111010000;
		weights[1200] <= 0000010100000000;
		weights[1201] <= 1000001010111011;
		weights[1202] <= 1000111111110111;
		weights[1203] <= 0000101110001011;
		weights[1204] <= 0001001111010000;
		weights[1205] <= 1001010101101011;
		weights[1206] <= 1000000101101011;
		weights[1207] <= 0000010001111011;
		weights[1208] <= 0000101001000101;
		weights[1209] <= 0000100000100101;
		weights[1210] <= 0000011110011110;
		weights[1211] <= 1000010010101010;
		weights[1212] <= 1000010011010101;
		weights[1213] <= 1000011100111011;
		weights[1214] <= 0000000101011000;
		weights[1215] <= 1000000111000001;
		weights[1216] <= 1000110101001001;
		weights[1217] <= 0000001111000111;
		weights[1218] <= 1000000000011110;
		weights[1219] <= 0000100100011001;
		weights[1220] <= 0000110111010011;
		weights[1221] <= 0000011000110000;
		weights[1222] <= 0000011101001001;
		weights[1223] <= 1000001111011101;
		weights[1224] <= 0000111001001101;
		weights[1225] <= 0000110000000100;
		weights[1226] <= 0000100000010000;
		weights[1227] <= 0000001110111101;
		weights[1228] <= 1000010000111011;
		weights[1229] <= 1000001110101000;
		weights[1230] <= 1000100001011011;
		weights[1231] <= 1000001100110110;
		weights[1232] <= 0000001110010111;
		weights[1233] <= 1000000011011100;
		weights[1234] <= 1000100001010000;
		weights[1235] <= 1000011001111010;
		weights[1236] <= 1000010001001101;
		weights[1237] <= 1000100010110110;
		weights[1238] <= 1000100100101100;
		weights[1239] <= 0000100111100000;
		weights[1240] <= 1000011010110110;
		weights[1241] <= 1000100001111101;
		weights[1242] <= 1000000001111000;
		weights[1243] <= 1000011011110110;
		weights[1244] <= 0001011101111101;
		weights[1245] <= 0000000111011011;
		weights[1246] <= 0000001001100110;
		weights[1247] <= 1000111001001100;
		weights[1248] <= 1000000000111010;
		weights[1249] <= 0000110101011100;
		weights[1250] <= 1000101001011111;
		weights[1251] <= 1000010110101100;
		weights[1252] <= 0000010110111110;
		weights[1253] <= 0000101110111111;
		weights[1254] <= 0000000100111010;
		weights[1255] <= 0000001001000111;
		weights[1256] <= 1000001011000010;
		weights[1257] <= 1000001110010000;
		weights[1258] <= 1000100011000100;
		weights[1259] <= 0000010110111111;
		weights[1260] <= 0001001001110100;
		weights[1261] <= 1001001100001001;
		weights[1262] <= 0000010011110100;
		weights[1263] <= 0000100011110000;
		weights[1264] <= 1001000111110100;
		weights[1265] <= 0000010001100000;
		weights[1266] <= 0000100101101101;
		weights[1267] <= 0000010000101101;
		weights[1268] <= 0000001110111010;
		weights[1269] <= 0000000010001011;
		weights[1270] <= 1000001011110010;
		weights[1271] <= 0000011101001110;
		weights[1272] <= 0000000000000010;
		weights[1273] <= 0000010101010010;
		weights[1274] <= 1000000110010000;
		weights[1275] <= 1000100010001100;
		weights[1276] <= 1000011011111111;
		weights[1277] <= 1000000111111110;
		weights[1278] <= 0000011110000100;
		weights[1279] <= 0000000010000011;
		weights[1280] <= 1000010111011110;
		weights[1281] <= 1000101011100110;
		weights[1282] <= 1000101110101100;
		weights[1283] <= 0000001010101101;
		weights[1284] <= 1000001110010110;
		weights[1285] <= 0000001101100110;
		weights[1286] <= 1000011111000101;
		weights[1287] <= 0000000111110000;
		weights[1288] <= 1000001100111101;
		weights[1289] <= 0000010001001010;
		weights[1290] <= 0001000001010110;
		weights[1291] <= 0000110111000000;
		weights[1292] <= 0000000100000110;
		weights[1293] <= 1000010001110100;
		weights[1294] <= 1000000111111011;
		weights[1295] <= 0000011000001111;
		weights[1296] <= 1000000010100100;
		weights[1297] <= 1000001110010111;
		weights[1298] <= 1000010110101000;
		weights[1299] <= 0001001011100011;
		weights[1300] <= 1000010111000000;
		weights[1301] <= 1000010011110010;
		weights[1302] <= 1000011001010110;
		weights[1303] <= 1000001000001001;
		weights[1304] <= 1000001001110100;
		weights[1305] <= 0000110001011001;
		weights[1306] <= 1000110001010001;
		weights[1307] <= 1000010010111110;
		weights[1308] <= 0000000101011111;
		weights[1309] <= 0000100001100000;
		weights[1310] <= 0000010000010011;
		weights[1311] <= 1000001001110111;
		weights[1312] <= 1000111101110000;
		weights[1313] <= 0000110000111111;
		weights[1314] <= 0000011100011000;
		weights[1315] <= 0000000110101100;
		weights[1316] <= 1000110011001111;
		weights[1317] <= 0000010100000101;
		weights[1318] <= 1000010110110111;
		weights[1319] <= 1000010111100010;
		weights[1320] <= 1000110000011101;
		weights[1321] <= 0000000001011100;
		weights[1322] <= 1000011000000000;
		weights[1323] <= 1000010111001101;
		weights[1324] <= 1000001110010111;
		weights[1325] <= 1000010001100011;
		weights[1326] <= 0000100110100101;
		weights[1327] <= 0000000010000000;
		weights[1328] <= 1000011010111011;
		weights[1329] <= 1000000000111001;
		weights[1330] <= 1000100010100101;
		weights[1331] <= 1000000010110010;
		weights[1332] <= 0000000010101010;
		weights[1333] <= 1000001000000001;
		weights[1334] <= 0000011001101000;
		weights[1335] <= 1000000110010001;
		weights[1336] <= 1000001001100001;
		weights[1337] <= 1000010111111011;
		weights[1338] <= 1000101000010101;
		weights[1339] <= 0000001000001000;
		weights[1340] <= 0000110011100001;
		weights[1341] <= 1000001101100100;
		weights[1342] <= 0000010111010101;
		weights[1343] <= 1000001100100100;
		weights[1344] <= 1000100100001100;
		weights[1345] <= 1000001100110111;
		weights[1346] <= 1000111111010011;
		weights[1347] <= 0000010001000101;
		weights[1348] <= 1000111011010000;
		weights[1349] <= 1000000010111000;
		weights[1350] <= 0000001111101011;
		weights[1351] <= 0000010001111100;
		weights[1352] <= 1001000101110100;
		weights[1353] <= 0000111000011011;
		weights[1354] <= 0000100011111110;
		weights[1355] <= 0000001101001001;
		weights[1356] <= 0000001100110111;
		weights[1357] <= 1000010101011100;
		weights[1358] <= 0000010101000000;
		weights[1359] <= 1000011100110100;
		weights[1360] <= 0000110111010011;
		weights[1361] <= 1000100001111010;
		weights[1362] <= 0000000100100101;
		weights[1363] <= 1000000000001011;
		weights[1364] <= 1000011001101100;
		weights[1365] <= 0000011001100001;
		weights[1366] <= 0000000111000000;
		weights[1367] <= 0000001101101011;
		weights[1368] <= 1000011001101001;
		weights[1369] <= 0000001001111010;
		weights[1370] <= 0000011000110101;
		weights[1371] <= 0000101100110101;
		weights[1372] <= 1000011110000001;
		weights[1373] <= 0000110010010101;
		weights[1374] <= 0000001100111111;
		weights[1375] <= 1000101000111100;
		weights[1376] <= 1000001100010000;
		weights[1377] <= 1000000110110101;
		weights[1378] <= 0000001001001011;
		weights[1379] <= 0000001011001010;
		weights[1380] <= 0001000100001100;
		weights[1381] <= 0000000001101110;
		weights[1382] <= 0000011000011101;
		weights[1383] <= 0000101000011101;
		weights[1384] <= 0000010000010101;
		weights[1385] <= 1000011110101111;
		weights[1386] <= 0000000111010010;
		weights[1387] <= 1000001001110111;
		weights[1388] <= 0000001011010011;
		weights[1389] <= 1000001010111010;
		weights[1390] <= 1000100010101111;
		weights[1391] <= 0000001100101110;
		weights[1392] <= 0000011011111100;
		weights[1393] <= 0000001100010110;
		weights[1394] <= 0000000010110111;
		weights[1395] <= 1000101100010110;
		weights[1396] <= 0000010011000110;
		weights[1397] <= 1000110101001100;
		weights[1398] <= 0000001100000100;
		weights[1399] <= 1000000110011101;
		weights[1400] <= 1000011011111010;
		weights[1401] <= 1000101111000010;
		weights[1402] <= 1000001001011001;
		weights[1403] <= 1000011011001011;
		weights[1404] <= 0000100011111010;
		weights[1405] <= 0000011110010111;
		weights[1406] <= 1000011101001100;
		weights[1407] <= 1000000110110101;
		weights[1408] <= 0000011111100100;
		weights[1409] <= 1000011011110111;
		weights[1410] <= 0000000111000011;
		weights[1411] <= 1000001010100111;
		weights[1412] <= 0000100110011100;
		weights[1413] <= 0000001111001101;
		weights[1414] <= 0000000111110101;
		weights[1415] <= 0001000010000101;
		weights[1416] <= 1000100101000110;
		weights[1417] <= 0000010101001111;
		weights[1418] <= 1000011000000101;
		weights[1419] <= 0000010001111100;
		weights[1420] <= 1000011111010000;
		weights[1421] <= 1000000000110100;
		weights[1422] <= 0000001001100110;
		weights[1423] <= 1000100110101111;
		weights[1424] <= 0000100000011001;
		weights[1425] <= 0000000100111010;
		weights[1426] <= 0000010011000111;
		weights[1427] <= 0000010101000101;
		weights[1428] <= 0000000100010101;
		weights[1429] <= 0001000001100011;
		weights[1430] <= 1000001100100010;
		weights[1431] <= 0000011001010110;
		weights[1432] <= 0000001010000101;
		weights[1433] <= 0000011110110101;
		weights[1434] <= 1000000000011111;
		weights[1435] <= 0000100011111001;
		weights[1436] <= 1000010000010011;
		weights[1437] <= 1000011110100101;
		weights[1438] <= 1000101011001001;
		weights[1439] <= 1000101011101111;
		weights[1440] <= 1000001100010000;
		weights[1441] <= 0000001010000000;
		weights[1442] <= 0000010101011100;
		weights[1443] <= 0001110111101111;
		weights[1444] <= 1000000101111011;
		weights[1445] <= 1000100010101001;
		weights[1446] <= 1000111111000000;
		weights[1447] <= 1000010110100010;
		weights[1448] <= 0000100011110110;
		weights[1449] <= 1000011101100110;
		weights[1450] <= 0000010000011011;
		weights[1451] <= 0000000101100100;
		weights[1452] <= 0000011101110000;
		weights[1453] <= 0000100111111101;
		weights[1454] <= 0000101111000010;
		weights[1455] <= 1000000111001011;
		weights[1456] <= 0000100101010101;
		weights[1457] <= 1000010011100000;
		weights[1458] <= 0000110000100101;
		weights[1459] <= 0000000100110010;
		weights[1460] <= 0000001011000001;
		weights[1461] <= 0000011001011100;
		weights[1462] <= 0000001100000000;
		weights[1463] <= 1000101100100111;
		weights[1464] <= 1000110110100000;
		weights[1465] <= 0000001001100100;
		weights[1466] <= 0000010010000001;
		weights[1467] <= 1000000100110000;
		weights[1468] <= 1000001000010100;
		weights[1469] <= 1000001101000010;
		weights[1470] <= 0000001100100001;
		weights[1471] <= 1000000100101101;
		weights[1472] <= 0000101110110100;
		weights[1473] <= 1000000000011001;
		weights[1474] <= 0000000101011001;
		weights[1475] <= 1000000000010110;
		weights[1476] <= 0000001001011010;
		weights[1477] <= 0000000110101101;
		weights[1478] <= 0000111010101011;
		weights[1479] <= 1000011101111001;
		weights[1480] <= 0000100101011001;
		weights[1481] <= 0000001001010111;
		weights[1482] <= 1000001010110110;
		weights[1483] <= 1000101010100110;
		weights[1484] <= 1000111001000100;
		weights[1485] <= 1000000111010111;
		weights[1486] <= 0000001000000011;
		weights[1487] <= 0000111000100101;
		weights[1488] <= 1000101001110101;
		weights[1489] <= 0000001001100100;
		weights[1490] <= 1000000110011101;
		weights[1491] <= 0000101010100001;
		weights[1492] <= 0000010110000011;
		weights[1493] <= 1000000110100011;
		weights[1494] <= 0000100010100101;
		weights[1495] <= 0000000101001011;
		weights[1496] <= 1000011111101100;
		weights[1497] <= 1000100111110100;
		weights[1498] <= 0000010010001000;
		weights[1499] <= 1000010111011011;
		weights[1500] <= 0000010010111000;
		weights[1501] <= 0000101011111011;
		weights[1502] <= 0000011110001100;
		weights[1503] <= 0000000111111111;
		weights[1504] <= 1000010011111011;
		weights[1505] <= 1000110000111000;
		weights[1506] <= 1000100001110101;
		weights[1507] <= 1000000010001101;
		weights[1508] <= 0000001010010011;
		weights[1509] <= 0000000110000000;
		weights[1510] <= 0000111110001111;
		weights[1511] <= 1000000001100100;
		weights[1512] <= 0000010010111000;
		weights[1513] <= 1000101100011100;
		weights[1514] <= 1000000001110000;
		weights[1515] <= 1000100100000001;
		weights[1516] <= 1000100111011111;
		weights[1517] <= 0000010011000101;
		weights[1518] <= 0001001100111100;
		weights[1519] <= 0000101010101101;
		weights[1520] <= 0000101000100010;
		weights[1521] <= 0000110000010011;
		weights[1522] <= 0000000000111110;
		weights[1523] <= 1000001010011111;
		weights[1524] <= 0000000001101100;
		weights[1525] <= 1000011111011101;
		weights[1526] <= 1000011100111111;
		weights[1527] <= 0000010011100001;
		weights[1528] <= 0000011001000001;
		weights[1529] <= 0000110101110010;
		weights[1530] <= 0000000111001110;
		weights[1531] <= 0000100110100111;
		weights[1532] <= 0000001010111010;
		weights[1533] <= 1000100010110110;
		weights[1534] <= 1000010010001010;
		weights[1535] <= 1000001011010100;
		weights[1536] <= 1000010100110010;
		weights[1537] <= 0000011100111100;
		weights[1538] <= 0000011010001110;
		weights[1539] <= 0000110100000111;
		weights[1540] <= 1000001011011001;
		weights[1541] <= 0000110100110110;
		weights[1542] <= 1000100000010000;
		weights[1543] <= 0000011011101110;
		weights[1544] <= 1000010011110001;
		weights[1545] <= 1000100111101001;
		weights[1546] <= 1000010001110011;
		weights[1547] <= 0000000111011110;
		weights[1548] <= 0000000011010011;
		weights[1549] <= 0000000011111010;
		weights[1550] <= 1000100111010010;
		weights[1551] <= 1000010000101111;
		weights[1552] <= 1000100010000000;
		weights[1553] <= 1000000110101000;
		weights[1554] <= 0000000110000110;
		weights[1555] <= 1000110010000001;
		weights[1556] <= 1000110000101001;
		weights[1557] <= 0000011111100010;
		weights[1558] <= 0000001101001010;
		weights[1559] <= 1000010111000101;
		weights[1560] <= 0000011101110100;
		weights[1561] <= 1000001000100100;
		weights[1562] <= 0000000011001001;
		weights[1563] <= 1000010010100110;
		weights[1564] <= 1000001101111001;
		weights[1565] <= 0000011000010011;
		weights[1566] <= 0000010111101111;
		weights[1567] <= 0000000101101010;
		weights[1568] <= 0000001111111111;
		weights[1569] <= 1000001100001110;
		weights[1570] <= 1000100010000111;
		weights[1571] <= 1000010011110101;
		weights[1572] <= 0000111010000110;
		weights[1573] <= 0000111100101100;
		weights[1574] <= 0001010100110011;
		weights[1575] <= 0000001100110011;
		weights[1576] <= 0000010011100100;
		weights[1577] <= 0000011101011101;
		weights[1578] <= 1000000111001011;
		weights[1579] <= 1000110001101011;
		weights[1580] <= 0000101100100000;
		weights[1581] <= 0000010000001001;
		weights[1582] <= 1000100110100111;
		weights[1583] <= 1000010110001100;
		weights[1584] <= 0000011111111001;
		weights[1585] <= 1000101110000010;
		weights[1586] <= 0000100100011000;
		weights[1587] <= 0001010010101101;
		weights[1588] <= 0000010111010001;
		weights[1589] <= 1000000000011100;
		weights[1590] <= 0000001111100110;
		weights[1591] <= 0000000111111000;
		weights[1592] <= 0000010010000010;
		weights[1593] <= 0000010011100010;
		weights[1594] <= 0000011010111010;
		weights[1595] <= 1000000011011001;
		weights[1596] <= 1000100110101100;
		weights[1597] <= 1000011110000100;
		weights[1598] <= 0000000010100011;
		weights[1599] <= 1000000010100101;
		weights[1600] <= 0000011011110110;
		weights[1601] <= 0000011111000011;
		weights[1602] <= 1000001110001010;
		weights[1603] <= 0001001000011000;
		weights[1604] <= 1000100010101010;
		weights[1605] <= 1000001101101100;
		weights[1606] <= 1000100001101110;
		weights[1607] <= 1000011100001101;
		weights[1608] <= 0000010110000100;
		weights[1609] <= 0000100100001101;
		weights[1610] <= 0000011000010000;
		weights[1611] <= 0000000010000000;
		weights[1612] <= 0000010001001000;
		weights[1613] <= 0000110010001010;
		weights[1614] <= 1000001101001110;
		weights[1615] <= 1001000000010100;
		weights[1616] <= 1000001101111101;
		weights[1617] <= 0000001101110011;
		weights[1618] <= 1000110010000000;
		weights[1619] <= 0000100011100101;
		weights[1620] <= 1000100000111111;
		weights[1621] <= 0000100001001001;
		weights[1622] <= 1000010010101100;
		weights[1623] <= 0000010100110100;
		weights[1624] <= 1000100001111010;
		weights[1625] <= 1000011111000001;
		weights[1626] <= 0000000011111101;
		weights[1627] <= 1000011101110110;
		weights[1628] <= 1000100010111110;
		weights[1629] <= 1000110101101101;
		weights[1630] <= 0000011110011110;
		weights[1631] <= 1000100000001011;
		weights[1632] <= 1000001011101011;
		weights[1633] <= 1000010100101001;
		weights[1634] <= 1000000111101010;
		weights[1635] <= 0000101111100011;
		weights[1636] <= 1001000001000111;
		weights[1637] <= 0000100111101101;
		weights[1638] <= 0000000111011000;
		weights[1639] <= 0000000011010010;
		weights[1640] <= 0000001111001001;
		weights[1641] <= 0000110110010100;
		weights[1642] <= 0000010011110110;
		weights[1643] <= 0000001101111101;
		weights[1644] <= 0000000101010101;
		weights[1645] <= 1000001010011011;
		weights[1646] <= 0000000011010100;
		weights[1647] <= 1000000101110111;
		weights[1648] <= 1000100111011111;
		weights[1649] <= 0000011001001101;
		weights[1650] <= 0000011110100101;
		weights[1651] <= 0000111000111010;
		weights[1652] <= 1000010101001011;
		weights[1653] <= 0000001110110111;
		weights[1654] <= 1000110010010101;
		weights[1655] <= 0000010110111010;
		weights[1656] <= 0000010001001001;
		weights[1657] <= 1000001111110010;
		weights[1658] <= 0000000101011101;
		weights[1659] <= 0000011100000010;
		weights[1660] <= 0000000010101100;
		weights[1661] <= 1000011001000000;
		weights[1662] <= 0000010101000100;
		weights[1663] <= 0000000011101000;
		weights[1664] <= 0000110100011010;
		weights[1665] <= 1000010001110000;
		weights[1666] <= 0000001001101111;
		weights[1667] <= 0000011010111011;
		weights[1668] <= 0000010110100010;
		weights[1669] <= 0000100100111101;
		weights[1670] <= 1000101000111001;
		weights[1671] <= 0000000100011101;
		weights[1672] <= 1000001001010110;
		weights[1673] <= 0000111100110001;
		weights[1674] <= 0000000001100001;
		weights[1675] <= 1000101010100001;
		weights[1676] <= 0000001010010000;
		weights[1677] <= 0000110011110010;
		weights[1678] <= 0000010011100001;
		weights[1679] <= 0001001100010110;
		weights[1680] <= 1000000101110111;
		weights[1681] <= 1000101110101110;
		weights[1682] <= 0000000111010011;
		weights[1683] <= 0000000010100010;
		weights[1684] <= 0000011000001111;
		weights[1685] <= 0000010011110100;
		weights[1686] <= 0000001011000111;
		weights[1687] <= 0000110110111010;
		weights[1688] <= 0000000111101111;
		weights[1689] <= 1000011100101001;
		weights[1690] <= 0000111001101111;
		weights[1691] <= 1000000110010101;
		weights[1692] <= 0000000000100011;
		weights[1693] <= 0001000110111110;
		weights[1694] <= 1000000010001100;
		weights[1695] <= 0000011011011110;
		weights[1696] <= 1000011010110000;
		weights[1697] <= 1000111001011010;
		weights[1698] <= 1000010010100001;
		weights[1699] <= 1000001100011001;
		weights[1700] <= 0000000100111110;
		weights[1701] <= 1000001001011100;
		weights[1702] <= 0000000111110101;
		weights[1703] <= 0000011110101110;
		weights[1704] <= 0000011100111011;
		weights[1705] <= 0000100010110011;
		weights[1706] <= 1000001011100000;
		weights[1707] <= 1000101011111110;
		weights[1708] <= 0000011110000110;
		weights[1709] <= 0000011100101011;
		weights[1710] <= 1000010011111010;
		weights[1711] <= 0000011101110111;
		weights[1712] <= 0000001110011000;
		weights[1713] <= 1000000100011011;
		weights[1714] <= 0000001101001110;
		weights[1715] <= 1000001101011011;
		weights[1716] <= 0000011011011011;
		weights[1717] <= 1000000011100110;
		weights[1718] <= 1000010110011010;
		weights[1719] <= 0000000100100110;
		weights[1720] <= 0000001000001111;
		weights[1721] <= 0000010111001000;
		weights[1722] <= 0000100000011000;
		weights[1723] <= 0000001001110011;
		weights[1724] <= 1000011100110110;
		weights[1725] <= 0000011110010011;
		weights[1726] <= 1000000011100011;
		weights[1727] <= 1000010010100011;
		weights[1728] <= 1000000011000101;
		weights[1729] <= 0000011101111000;
		weights[1730] <= 0000010011010000;
		weights[1731] <= 0000011001011100;
		weights[1732] <= 0000010000000110;
		weights[1733] <= 0000000101111010;
		weights[1734] <= 1000001100111010;
		weights[1735] <= 1000000011011110;
		weights[1736] <= 0000000000010100;
		weights[1737] <= 0000001011111110;
		weights[1738] <= 1000000011111011;
		weights[1739] <= 0000010001001110;
		weights[1740] <= 1000101101111100;
		weights[1741] <= 1000001101101011;
		weights[1742] <= 0000100000011100;
		weights[1743] <= 0000010101101101;
		weights[1744] <= 1000011111010000;
		weights[1745] <= 1001100101001001;
		weights[1746] <= 0000010101000011;
		weights[1747] <= 0000101100110110;
		weights[1748] <= 0000010010010010;
		weights[1749] <= 0000010000010101;
		weights[1750] <= 0000010001011001;
		weights[1751] <= 0000011010011001;
		weights[1752] <= 0000000010000100;
		weights[1753] <= 1000000011111111;
		weights[1754] <= 1000001000000011;
		weights[1755] <= 1000000001100001;
		weights[1756] <= 1000001000011101;
		weights[1757] <= 1000001111001011;
		weights[1758] <= 0000000100000001;
		weights[1759] <= 0000000100101111;
		weights[1760] <= 0001000101110010;
		weights[1761] <= 0000100110000100;
		weights[1762] <= 1000001110010111;
		weights[1763] <= 0001010001100010;
		weights[1764] <= 1000001010110000;
		weights[1765] <= 1000011000101101;
		weights[1766] <= 1000001001101011;
		weights[1767] <= 1000000101100001;
		weights[1768] <= 0000100101111111;
		weights[1769] <= 0000000101011101;
		weights[1770] <= 0000001110000111;
		weights[1771] <= 0000001010010010;
		weights[1772] <= 0000101000001100;
		weights[1773] <= 0000001100110110;
		weights[1774] <= 0000011111001101;
		weights[1775] <= 0000000111010010;
		weights[1776] <= 0000101010001000;
		weights[1777] <= 0000100100110110;
		weights[1778] <= 0000010011101110;
		weights[1779] <= 1000111001101101;
		weights[1780] <= 1000110111110011;
		weights[1781] <= 1000011101011001;
		weights[1782] <= 1000000100010001;
		weights[1783] <= 1000011101011101;
		weights[1784] <= 0000010011001110;
		weights[1785] <= 0000110100010110;
		weights[1786] <= 0000001100000111;
		weights[1787] <= 1000010101000110;
		weights[1788] <= 0000011001000111;
		weights[1789] <= 1000001000110011;
		weights[1790] <= 1000000110111011;
		weights[1791] <= 0000001110010011;
		weights[1792] <= 0000100100001101;
		weights[1793] <= 0001010010111001;
		weights[1794] <= 0001001110011110;
		weights[1795] <= 0001011101110000;
		weights[1796] <= 0001010111000101;
		weights[1797] <= 1000100111010111;
		weights[1798] <= 0000000110100110;
		weights[1799] <= 1000010001100111;
		weights[1800] <= 0001000011001010;
		weights[1801] <= 0000001110000000;
		weights[1802] <= 0000000001111001;
		weights[1803] <= 0000101100111110;
		weights[1804] <= 1000000011110001;
		weights[1805] <= 0000101000010111;
		weights[1806] <= 0000001111110001;
		weights[1807] <= 1000000000001010;
		weights[1808] <= 1000010000111110;
		weights[1809] <= 1000010001010001;
		weights[1810] <= 1000110010111010;
		weights[1811] <= 1000000001110101;
		weights[1812] <= 0000000010111110;
		weights[1813] <= 0001011010101001;
		weights[1814] <= 0000111010000110;
		weights[1815] <= 0001010111101000;
		weights[1816] <= 1000010101000011;
		weights[1817] <= 1000000000000100;
		weights[1818] <= 0000010000011010;
		weights[1819] <= 1000010001110011;
		weights[1820] <= 0000011010010010;
		weights[1821] <= 0000101011000000;
		weights[1822] <= 1000000011000011;
		weights[1823] <= 0001011011111101;
		weights[1824] <= 1000001000110001;
		weights[1825] <= 1000101001011101;
		weights[1826] <= 0000000111110000;
		weights[1827] <= 0000010000001111;
		weights[1828] <= 0000001011011000;
		weights[1829] <= 1000011000011110;
		weights[1830] <= 1000001111001010;
		weights[1831] <= 1000001110100111;
		weights[1832] <= 0000000001001001;
		weights[1833] <= 0000000110001011;
		weights[1834] <= 0000010010110001;
		weights[1835] <= 0000011111110010;
		weights[1836] <= 0000010000011001;
		weights[1837] <= 1000000010011101;
		weights[1838] <= 0000000010000100;
		weights[1839] <= 1000001011100111;
		weights[1840] <= 1000010101111000;
		weights[1841] <= 0000000110110010;
		weights[1842] <= 1000101111100110;
		weights[1843] <= 1000010111100010;
		weights[1844] <= 0000010001100010;
		weights[1845] <= 0000010010000101;
		weights[1846] <= 1000010001111011;
		weights[1847] <= 1000100110011101;
		weights[1848] <= 1000001100101000;
		weights[1849] <= 1000010101101010;
		weights[1850] <= 1000001010110001;
		weights[1851] <= 1000000001011111;
		weights[1852] <= 1000001010011101;
		weights[1853] <= 1000011000100011;
		weights[1854] <= 0000010111111110;
		weights[1855] <= 0000000010001001;
		weights[1856] <= 0000001001000101;
		weights[1857] <= 0000000010010110;
		weights[1858] <= 0000001000010010;
		weights[1859] <= 0000000010010010;
		weights[1860] <= 1000100100011011;
		weights[1861] <= 1000001101010010;
		weights[1862] <= 0000010111011011;
		weights[1863] <= 0000100111011100;
		weights[1864] <= 0000001000010100;
		weights[1865] <= 0000001011110001;
		weights[1866] <= 1000000001111100;
		weights[1867] <= 0000011110110101;
		weights[1868] <= 1000001111100111;
		weights[1869] <= 1000001011101111;
		weights[1870] <= 0000000011100111;
		weights[1871] <= 0000010111011101;
		weights[1872] <= 0000001001010001;
		weights[1873] <= 1000010010111111;
		weights[1874] <= 0000000010111100;
		weights[1875] <= 1000001010100010;
		weights[1876] <= 0000001000010111;
		weights[1877] <= 1000001011111110;
		weights[1878] <= 0000000111001110;
		weights[1879] <= 0000001001101000;
		weights[1880] <= 0000101001000000;
		weights[1881] <= 0000000110101011;
		weights[1882] <= 1000000010110100;
		weights[1883] <= 1000000110011011;
		weights[1884] <= 1000011110110101;
		weights[1885] <= 0000100110100111;
		weights[1886] <= 1000001110001011;
		weights[1887] <= 1000001001111111;
		weights[1888] <= 1000001101101101;
		weights[1889] <= 0000001011101100;
		weights[1890] <= 0000000111100010;
		weights[1891] <= 1000000101101011;
		weights[1892] <= 0000011111101001;
		weights[1893] <= 1000000010101011;
		weights[1894] <= 1000011100111110;
		weights[1895] <= 0000000011100100;
		weights[1896] <= 0000011000111000;
		weights[1897] <= 0000001001010000;
		weights[1898] <= 1000101100010100;
		weights[1899] <= 0000011111001010;
		weights[1900] <= 1000000111100001;
		weights[1901] <= 0000011011101101;
		weights[1902] <= 1000000000111010;
		weights[1903] <= 1001000001001011;
		weights[1904] <= 1000001011001101;
		weights[1905] <= 0000110010010110;
		weights[1906] <= 1000011110101001;
		weights[1907] <= 0000000110011000;
		weights[1908] <= 1000011010110100;
		weights[1909] <= 1000001111011101;
		weights[1910] <= 0000011011000100;
		weights[1911] <= 1000010000000111;
		weights[1912] <= 0000000001011000;
		weights[1913] <= 1000101001001001;
		weights[1914] <= 0000001110101000;
		weights[1915] <= 0000010110111000;
		weights[1916] <= 1000010000100011;
		weights[1917] <= 1000010011111001;
		weights[1918] <= 0000001101111001;
		weights[1919] <= 1000000111100100;
		weights[1920] <= 0000001100001011;
		weights[1921] <= 1000010101000111;
		weights[1922] <= 0000000011110101;
		weights[1923] <= 1000101001100001;
		weights[1924] <= 1000001010100111;
		weights[1925] <= 0000001001101001;
		weights[1926] <= 0000010001110011;
		weights[1927] <= 1000011010111000;
		weights[1928] <= 0000101101101000;
		weights[1929] <= 1000110011010111;
		weights[1930] <= 0001000111101000;
		weights[1931] <= 1000000101011010;
		weights[1932] <= 0000001101001010;
		weights[1933] <= 0000011001001011;
		weights[1934] <= 1000001100000001;
		weights[1935] <= 1000011111000101;
		weights[1936] <= 0000000011000010;
		weights[1937] <= 0000010001100001;
		weights[1938] <= 1000000100010000;
		weights[1939] <= 1000000010111001;
		weights[1940] <= 0000011010111101;
		weights[1941] <= 1000010100001100;
		weights[1942] <= 0000110100110111;
		weights[1943] <= 1000000001100011;
		weights[1944] <= 1000000100111011;
		weights[1945] <= 1000111100001001;
		weights[1946] <= 0000000001101010;
		weights[1947] <= 1000110001110101;
		weights[1948] <= 0000011010100010;
		weights[1949] <= 0000011011100010;
		weights[1950] <= 1000101100100001;
		weights[1951] <= 0000110100101011;
		weights[1952] <= 1000001000000111;
		weights[1953] <= 0000011011111110;
		weights[1954] <= 0000101110111010;
		weights[1955] <= 0000000111001100;
		weights[1956] <= 0000010000010000;
		weights[1957] <= 1000001001000000;
		weights[1958] <= 1000011110001011;
		weights[1959] <= 0001101101111110;
		weights[1960] <= 1000001000101011;
		weights[1961] <= 1000010011110100;
		weights[1962] <= 0000110100011010;
		weights[1963] <= 0000011110110010;
		weights[1964] <= 0000010100001010;
		weights[1965] <= 1000001011111010;
		weights[1966] <= 0000000111100100;
		weights[1967] <= 0000010111100111;
		weights[1968] <= 0000011101111001;
		weights[1969] <= 0000000000100101;
		weights[1970] <= 0001001110010001;
		weights[1971] <= 1000001110101101;
		weights[1972] <= 1000010001011100;
		weights[1973] <= 1000001100001011;
		weights[1974] <= 1000011001100100;
		weights[1975] <= 0000001011000101;
		weights[1976] <= 0000010101111100;
		weights[1977] <= 0000000000000001;
		weights[1978] <= 0001010100001010;
		weights[1979] <= 0001000100000011;
		weights[1980] <= 1000001111101100;
		weights[1981] <= 0000011001000010;
		weights[1982] <= 0001100101011100;
		weights[1983] <= 1000100011111011;
		weights[1984] <= 1000101011011101;
		weights[1985] <= 0000011110111011;
		weights[1986] <= 1000000111100001;
		weights[1987] <= 1000100000110101;
		weights[1988] <= 1000011100111011;
		weights[1989] <= 0000000011101000;
		weights[1990] <= 1000100111011001;
		weights[1991] <= 1000011001100100;
		weights[1992] <= 1000000010001110;
		weights[1993] <= 1000011010010000;
		weights[1994] <= 1000010100010001;
		weights[1995] <= 0000000011000101;
		weights[1996] <= 1000011110100000;
		weights[1997] <= 0000000101011011;
		weights[1998] <= 1000000001111000;
		weights[1999] <= 0000111010000000;
		weights[2000] <= 0000001011010110;
		weights[2001] <= 1000001100000101;
		weights[2002] <= 1000001010100011;
		weights[2003] <= 0000011011000111;
		weights[2004] <= 1010010011011000;
		weights[2005] <= 0000100011110000;
		weights[2006] <= 0000010010000101;
		weights[2007] <= 1000100100010100;
		weights[2008] <= 1000010100011011;
		weights[2009] <= 0000001100110110;
		weights[2010] <= 1000011000011001;
		weights[2011] <= 0000010001001110;
		weights[2012] <= 0000101110011110;
		weights[2013] <= 0000001101111000;
		weights[2014] <= 1000110000011110;
		weights[2015] <= 0001000111001101;
		weights[2016] <= 1001010100101111;
		weights[2017] <= 0000001010011111;
		weights[2018] <= 1000001101001101;
		weights[2019] <= 1000001101010000;
		weights[2020] <= 1000100011000001;
		weights[2021] <= 0000000001110001;
		weights[2022] <= 0000111110100110;
		weights[2023] <= 0000000110001110;
		weights[2024] <= 1000001110000101;
		weights[2025] <= 0000110001101010;
		weights[2026] <= 1000001001010111;
		weights[2027] <= 1000010101000011;
		weights[2028] <= 0000001110100010;
		weights[2029] <= 0000010110011111;
		weights[2030] <= 0000011111001011;
		weights[2031] <= 1000110100001100;
		weights[2032] <= 1000001101000101;
		weights[2033] <= 0000100000111000;
		weights[2034] <= 0000011101001100;
		weights[2035] <= 1000000100010101;
		weights[2036] <= 1000000011100001;
		weights[2037] <= 1000000101010101;
		weights[2038] <= 1000011010011100;
		weights[2039] <= 0000101000111111;
		weights[2040] <= 1000010110101111;
		weights[2041] <= 1000000110101111;
		weights[2042] <= 0000101000011010;
		weights[2043] <= 0000011001111111;
		weights[2044] <= 1000000111110000;
		weights[2045] <= 0000010000101101;
		weights[2046] <= 0000001100000111;
		weights[2047] <= 0001001001001110;
		weights[2048] <= 0000011001101101;
		weights[2049] <= 1000000100111101;
		weights[2050] <= 0000011000001100;
		weights[2051] <= 1000101011011001;
		weights[2052] <= 1000011101001110;
		weights[2053] <= 1000001011011100;
		weights[2054] <= 0000101001011100;
		weights[2055] <= 0000001000111110;
		weights[2056] <= 0000110010010001;
		weights[2057] <= 0000010110110001;
		weights[2058] <= 1000000101111101;
		weights[2059] <= 1000101011001110;
		weights[2060] <= 1000101100010100;
		weights[2061] <= 1000010101011000;
		weights[2062] <= 1000000001001011;
		weights[2063] <= 0000000001100101;
		weights[2064] <= 1000000001110111;
		weights[2065] <= 0000101100011001;
		weights[2066] <= 0000001111001110;
		weights[2067] <= 1000010101011100;
		weights[2068] <= 1000011001010011;
		weights[2069] <= 1000000101110001;
		weights[2070] <= 0000110100111101;
		weights[2071] <= 0000010110100011;
		weights[2072] <= 1000101010110010;
		weights[2073] <= 0000001000101101;
		weights[2074] <= 0000000001111000;
		weights[2075] <= 1000110001111100;
		weights[2076] <= 1000110111011010;
		weights[2077] <= 1000111110111010;
		weights[2078] <= 1000000011010101;
		weights[2079] <= 0000000010000111;
		weights[2080] <= 0000101110100110;
		weights[2081] <= 0000100110101111;
		weights[2082] <= 1000110001100110;
		weights[2083] <= 0000100110100111;
		weights[2084] <= 1000001101101001;
		weights[2085] <= 1000011011000001;
		weights[2086] <= 0000001101000001;
		weights[2087] <= 0000000010101010;
		weights[2088] <= 1000010000011001;
		weights[2089] <= 1000101100111010;
		weights[2090] <= 0000011011111101;
		weights[2091] <= 0000011001111110;
		weights[2092] <= 0000000001011100;
		weights[2093] <= 1000011101100110;
		weights[2094] <= 0000010111111000;
		weights[2095] <= 1000001001011011;
		weights[2096] <= 1000110101001011;
		weights[2097] <= 1000011000001010;
		weights[2098] <= 1000001100010000;
		weights[2099] <= 1000100110000001;
		weights[2100] <= 1000010111000011;
		weights[2101] <= 1000001101000001;
		weights[2102] <= 1000000111010001;
		weights[2103] <= 0000010000010100;
		weights[2104] <= 1000011000101011;
		weights[2105] <= 0000010001110011;
		weights[2106] <= 0000000011001001;
		weights[2107] <= 1000001110010001;
		weights[2108] <= 0000110011000001;
		weights[2109] <= 0000000010000000;
		weights[2110] <= 0000100101101100;
		weights[2111] <= 0000100001101011;
		weights[2112] <= 0000011001110011;
		weights[2113] <= 0000010110010110;
		weights[2114] <= 0000001010100101;
		weights[2115] <= 0000000011100101;
		weights[2116] <= 1000101101100011;
		weights[2117] <= 0000010111011010;
		weights[2118] <= 0000000000001101;
		weights[2119] <= 0000100010111100;
		weights[2120] <= 0000000100001010;
		weights[2121] <= 1000111100000000;
		weights[2122] <= 0000101101010000;
		weights[2123] <= 0000011100000110;
		weights[2124] <= 1000010100001101;
		weights[2125] <= 0000000101010010;
		weights[2126] <= 1000010101011001;
		weights[2127] <= 1000011010010001;
		weights[2128] <= 0000001010001000;
		weights[2129] <= 1000000111001100;
		weights[2130] <= 0000000011010011;
		weights[2131] <= 0000010010100000;
		weights[2132] <= 0000110101100011;
		weights[2133] <= 0000011110100000;
		weights[2134] <= 1000001010010111;
		weights[2135] <= 1000000100011000;
		weights[2136] <= 0000010001011000;
		weights[2137] <= 1000011000100001;
		weights[2138] <= 0000001000101001;
		weights[2139] <= 1000010010010111;
		weights[2140] <= 1000001110101001;
		weights[2141] <= 0000000001111000;
		weights[2142] <= 1000011110111110;
		weights[2143] <= 0000110000000001;
		weights[2144] <= 1000100000010101;
		weights[2145] <= 0000000010011110;
		weights[2146] <= 0000011111100010;
		weights[2147] <= 0000011011100111;
		weights[2148] <= 1000000011010110;
		weights[2149] <= 1000010000000101;
		weights[2150] <= 0000011001010010;
		weights[2151] <= 0000100101110000;
		weights[2152] <= 0000101001000100;
		weights[2153] <= 0000011110100101;
		weights[2154] <= 0000011101010111;
		weights[2155] <= 0000001011010110;
		weights[2156] <= 1000011101010011;
		weights[2157] <= 1000001111101011;
		weights[2158] <= 1000111111011011;
		weights[2159] <= 0000011100101001;
		weights[2160] <= 0000000110111110;
		weights[2161] <= 1000010101111101;
		weights[2162] <= 1000000101010111;
		weights[2163] <= 1000110001101000;
		weights[2164] <= 0000000110001100;
		weights[2165] <= 1000011011000001;
		weights[2166] <= 0000100101111110;
		weights[2167] <= 1000000000001101;
		weights[2168] <= 0000110001010001;
		weights[2169] <= 0000101101110011;
		weights[2170] <= 0000010000000111;
		weights[2171] <= 0000000010001011;
		weights[2172] <= 1000101001000010;
		weights[2173] <= 1000001001010010;
		weights[2174] <= 0000011111100111;
		weights[2175] <= 0000001011110100;
		weights[2176] <= 1001100101010011;
		weights[2177] <= 1000101101100101;
		weights[2178] <= 1000001101100101;
		weights[2179] <= 0000001100001000;
		weights[2180] <= 0000100000100010;
		weights[2181] <= 1000101100111010;
		weights[2182] <= 0000001000100110;
		weights[2183] <= 1000110100011001;
		weights[2184] <= 0000110000010110;
		weights[2185] <= 0000011101101110;
		weights[2186] <= 1000101101110011;
		weights[2187] <= 0000101100011010;
		weights[2188] <= 0000000011010110;
		weights[2189] <= 0000011010010101;
		weights[2190] <= 0000100100011110;
		weights[2191] <= 0000101010101000;
		weights[2192] <= 0000100111010100;
		weights[2193] <= 0000101010000011;
		weights[2194] <= 1000001101011111;
		weights[2195] <= 1000010011010111;
		weights[2196] <= 1000001000101111;
		weights[2197] <= 1000100111110011;
		weights[2198] <= 0000010110010110;
		weights[2199] <= 1000100010001100;
		weights[2200] <= 1001000010111111;
		weights[2201] <= 0000100101010000;
		weights[2202] <= 0000001010010001;
		weights[2203] <= 0000100111110111;
		weights[2204] <= 1000001110101010;
		weights[2205] <= 1000001110000001;
		weights[2206] <= 1000011101101100;
		weights[2207] <= 1000111001011100;
		weights[2208] <= 1000110000011101;
		weights[2209] <= 1000001011110000;
		weights[2210] <= 1000100001110011;
		weights[2211] <= 0000000100111011;
		weights[2212] <= 1000100100010011;
		weights[2213] <= 1000010110101111;
		weights[2214] <= 1000001101010110;
		weights[2215] <= 1000000101001011;
		weights[2216] <= 1000110100110010;
		weights[2217] <= 1000100101100100;
		weights[2218] <= 1000000000011111;
		weights[2219] <= 0000011001101011;
		weights[2220] <= 1000000101110000;
		weights[2221] <= 1000000010010001;
		weights[2222] <= 1000111001110111;
		weights[2223] <= 0000011010001001;
		weights[2224] <= 0000101001000111;
		weights[2225] <= 0000111010110010;
		weights[2226] <= 1000011011111010;
		weights[2227] <= 0000011110100101;
		weights[2228] <= 0000010110001011;
		weights[2229] <= 0000010001101001;
		weights[2230] <= 0000011010010000;
		weights[2231] <= 1000011000111010;
		weights[2232] <= 0000100110100100;
		weights[2233] <= 1000100011010111;
		weights[2234] <= 0000001011010101;
		weights[2235] <= 0000000000010000;
		weights[2236] <= 0000010000101001;
		weights[2237] <= 0000011001010110;
		weights[2238] <= 0000111100101101;
		weights[2239] <= 0000011001001000;
		weights[2240] <= 1000110010011001;
		weights[2241] <= 1000011010101110;
		weights[2242] <= 0000101010111101;
		weights[2243] <= 0000000010101010;
		weights[2244] <= 0000010001100110;
		weights[2245] <= 0000010111000100;
		weights[2246] <= 1000010000111010;
		weights[2247] <= 1000001110111000;
		weights[2248] <= 0000010100000000;
		weights[2249] <= 1000000100010000;
		weights[2250] <= 1000011111101101;
		weights[2251] <= 0000000100010000;
		weights[2252] <= 1000001111000011;
		weights[2253] <= 1000000001111001;
		weights[2254] <= 0000001010001111;
		weights[2255] <= 0000010011001010;
		weights[2256] <= 0000001011110011;
		weights[2257] <= 0000100101110010;
		weights[2258] <= 1000001110001001;
		weights[2259] <= 1001001101111100;
		weights[2260] <= 1000011011100011;
		weights[2261] <= 0000001100110011;
		weights[2262] <= 1000100101001000;
		weights[2263] <= 0000011000000000;
		weights[2264] <= 0000010010100101;
		weights[2265] <= 0000100011110000;
		weights[2266] <= 0000011010110010;
		weights[2267] <= 1000000101100101;
		weights[2268] <= 1000001001000110;
		weights[2269] <= 0000101101110100;
		weights[2270] <= 1000010011100101;
		weights[2271] <= 1000000101001000;
		weights[2272] <= 1000000100001001;
		weights[2273] <= 0000110000000011;
		weights[2274] <= 1000010101011001;
		weights[2275] <= 1000001010000001;
		weights[2276] <= 1000001011000011;
		weights[2277] <= 1000001010010011;
		weights[2278] <= 1000010100110011;
		weights[2279] <= 1000000111010111;
		weights[2280] <= 1000011101000100;
		weights[2281] <= 1000100001100000;
		weights[2282] <= 1000010110011000;
		weights[2283] <= 1000000110110011;
		weights[2284] <= 0000100101100110;
		weights[2285] <= 1001010111001000;
		weights[2286] <= 0000010100110110;
		weights[2287] <= 0000000111010000;
		weights[2288] <= 1000101011000110;
		weights[2289] <= 1000000001011011;
		weights[2290] <= 1000101101101010;
		weights[2291] <= 1000000111101000;
		weights[2292] <= 0000110101000010;
		weights[2293] <= 0000000001001110;
		weights[2294] <= 1000010000000110;
		weights[2295] <= 0000010110011100;
		weights[2296] <= 1000001110110110;
		weights[2297] <= 1000000100111010;
		weights[2298] <= 1000100010010011;
		weights[2299] <= 0000101110101101;
		weights[2300] <= 0000010110100001;
		weights[2301] <= 0000111010011001;
		weights[2302] <= 0000001100111101;
		weights[2303] <= 0000010110000111;
		weights[2304] <= 1000000101100110;
		weights[2305] <= 0001001000000111;
		weights[2306] <= 1000001010111011;
		weights[2307] <= 0000001010110001;
		weights[2308] <= 1000101110010001;
		weights[2309] <= 1000000010111010;
		weights[2310] <= 1000100010110100;
		weights[2311] <= 0000111111101101;
		weights[2312] <= 1000010000000010;
		weights[2313] <= 0001001001100001;
		weights[2314] <= 0000010000001111;
		weights[2315] <= 0000001000111010;
		weights[2316] <= 1000111111001011;
		weights[2317] <= 1000111010100011;
		weights[2318] <= 1000001011101101;
		weights[2319] <= 1000100001000111;
		weights[2320] <= 0000101111110101;
		weights[2321] <= 1000010001000111;
		weights[2322] <= 1000010101001001;
		weights[2323] <= 0000000100010010;
		weights[2324] <= 1000000100101010;
		weights[2325] <= 0000011001110011;
		weights[2326] <= 1000110111000100;
		weights[2327] <= 1000101101111000;
		weights[2328] <= 1000001001110001;
		weights[2329] <= 0000000001001111;
		weights[2330] <= 0000101011000101;
		weights[2331] <= 1000000100011100;
		weights[2332] <= 0000011011111000;
		weights[2333] <= 1000000111001000;
		weights[2334] <= 0000011101001010;
		weights[2335] <= 0000100110000101;
		weights[2336] <= 1000001011111001;
		weights[2337] <= 0000011000010011;
		weights[2338] <= 0000000101010000;
		weights[2339] <= 1000010010100110;
		weights[2340] <= 1000010000101101;
		weights[2341] <= 0000000111001000;
		weights[2342] <= 1000001111110101;
		weights[2343] <= 1000101101111001;
		weights[2344] <= 1001001100110001;
		weights[2345] <= 1000001111101011;
		weights[2346] <= 1000010100011101;
		weights[2347] <= 0000011101000101;
		weights[2348] <= 1000001100111011;
		weights[2349] <= 1000001101011001;
		weights[2350] <= 1000011101101000;
		weights[2351] <= 0000000110100110;
		weights[2352] <= 1000011110001101;
		weights[2353] <= 1000001010100010;
		weights[2354] <= 0000001100100111;
		weights[2355] <= 0000011101001011;
		weights[2356] <= 0000100110001000;
		weights[2357] <= 0000010100011111;
		weights[2358] <= 0000001001010111;
		weights[2359] <= 0000011110110111;
		weights[2360] <= 1000010100011110;
		weights[2361] <= 0000000111111100;
		weights[2362] <= 0000111010001100;
		weights[2363] <= 1000010110011111;
		weights[2364] <= 0000001001000111;
		weights[2365] <= 0000001000011100;
		weights[2366] <= 0000000110000010;
		weights[2367] <= 1000110110101100;
		weights[2368] <= 1000011100011101;
		weights[2369] <= 1000010101110101;
		weights[2370] <= 1000110010100110;
		weights[2371] <= 1000100111010101;
		weights[2372] <= 0000100000000011;
		weights[2373] <= 1000100101010100;
		weights[2374] <= 0000011001011110;
		weights[2375] <= 1000110101111110;
		weights[2376] <= 0000001101101000;
		weights[2377] <= 0000110100011011;
		weights[2378] <= 0000010101101011;
		weights[2379] <= 1000010111100111;
		weights[2380] <= 1000011101101101;
		weights[2381] <= 0000001001100000;
		weights[2382] <= 1000011000001011;
		weights[2383] <= 1000100101011000;
		weights[2384] <= 0000011101000000;
		weights[2385] <= 1000000010110111;
		weights[2386] <= 0000010001111110;
		weights[2387] <= 1000000100100000;
		weights[2388] <= 0001001000001110;
		weights[2389] <= 0000001011111000;
		weights[2390] <= 1000001010001010;
		weights[2391] <= 0000100000011001;
		weights[2392] <= 1000000000110011;
		weights[2393] <= 1000001110000010;
		weights[2394] <= 1000000111000000;
		weights[2395] <= 1000010000000110;
		weights[2396] <= 1000111110101011;
		weights[2397] <= 1000100000001000;
		weights[2398] <= 1000001100111010;
		weights[2399] <= 0000000110111011;
		weights[2400] <= 1000001100110000;
		weights[2401] <= 1000101001101110;
		weights[2402] <= 1000001011100001;
		weights[2403] <= 1000001101011011;
		weights[2404] <= 0000000000100100;
		weights[2405] <= 0001001001011000;
		weights[2406] <= 0000000101010110;
		weights[2407] <= 1000000001011101;
		weights[2408] <= 0000100011011110;
		weights[2409] <= 1000000100011000;
		weights[2410] <= 0000011000011011;
		weights[2411] <= 1000000011010010;
		weights[2412] <= 0000011100110011;
		weights[2413] <= 0000001101100110;
		weights[2414] <= 1000001001000111;
		weights[2415] <= 1000001110110010;
		weights[2416] <= 0000001000011001;
		weights[2417] <= 0000001100111110;
		weights[2418] <= 0000000100101110;
		weights[2419] <= 1000001100110011;
		weights[2420] <= 0001001110111100;
		weights[2421] <= 1000000101110111;
		weights[2422] <= 0000101101111110;
		weights[2423] <= 0000010110001101;
		weights[2424] <= 0000001011111001;
		weights[2425] <= 0000111110100100;
		weights[2426] <= 1000111001111010;
		weights[2427] <= 1000000100111101;
		weights[2428] <= 0000110000011101;
		weights[2429] <= 1000001101001000;
		weights[2430] <= 0000111100000100;
		weights[2431] <= 1000101100001110;
		weights[2432] <= 1000001111110010;
		weights[2433] <= 0000011100010110;
		weights[2434] <= 0000011100011011;
		weights[2435] <= 0000001000110101;
		weights[2436] <= 0000011100110001;
		weights[2437] <= 0000001000010000;
		weights[2438] <= 0000010100101000;
		weights[2439] <= 1000101101101100;
		weights[2440] <= 0000001011010100;
		weights[2441] <= 1000010101100010;
		weights[2442] <= 0000001001010000;
		weights[2443] <= 0000101110011000;
		weights[2444] <= 0000001100101000;
		weights[2445] <= 0000000101110101;
		weights[2446] <= 0000011001101000;
		weights[2447] <= 0000100010000110;
		weights[2448] <= 1000001100111100;
		weights[2449] <= 0000110000010101;
		weights[2450] <= 0000001100001110;
		weights[2451] <= 1000100010010000;
		weights[2452] <= 1000010101000110;
		weights[2453] <= 0000010000110110;
		weights[2454] <= 1000011000111001;
		weights[2455] <= 1000100100100011;
		weights[2456] <= 1000000100001101;
		weights[2457] <= 0000110101111110;
		weights[2458] <= 0000001110100001;
		weights[2459] <= 1000000010111110;
		weights[2460] <= 0000110001111101;
		weights[2461] <= 1000011111101001;
		weights[2462] <= 1000101100000111;
		weights[2463] <= 1001000000010011;
		weights[2464] <= 0000000111111011;
		weights[2465] <= 1000010110011101;
		weights[2466] <= 0000011111001110;
		weights[2467] <= 0000001111011100;
		weights[2468] <= 0000010110110011;
		weights[2469] <= 1000001000001101;
		weights[2470] <= 0000000110000101;
		weights[2471] <= 1000101110100010;
		weights[2472] <= 0000100101011100;
		weights[2473] <= 1000000111010101;
		weights[2474] <= 0000100011010111;
		weights[2475] <= 1000001100110010;
		weights[2476] <= 1000100110011001;
		weights[2477] <= 1000010101111111;
		weights[2478] <= 0000011011010110;
		weights[2479] <= 0000010001000110;
		weights[2480] <= 1000010100000111;
		weights[2481] <= 0000000101001110;
		weights[2482] <= 1000000101000101;
		weights[2483] <= 0000000000101011;
		weights[2484] <= 1000011010110101;
		weights[2485] <= 0000001001110101;
		weights[2486] <= 1000010100001111;
		weights[2487] <= 0000010010101101;
		weights[2488] <= 1000010011110101;
		weights[2489] <= 0000000011101000;
		weights[2490] <= 1000101111011000;
		weights[2491] <= 1000101100011000;
		weights[2492] <= 1000101100100111;
		weights[2493] <= 1000001011111100;
		weights[2494] <= 0000110111111111;
		weights[2495] <= 0000001100000110;
		weights[2496] <= 1000010011010110;
		weights[2497] <= 1000110110100011;
		weights[2498] <= 1000010110000000;
		weights[2499] <= 1001001010011000;
		weights[2500] <= 1000101011101010;
		weights[2501] <= 1000000110000101;
		weights[2502] <= 0000101001110011;
		weights[2503] <= 0000100101110101;
		weights[2504] <= 0000110001000101;
		weights[2505] <= 0000010110001100;
		weights[2506] <= 0000010101001111;
		weights[2507] <= 1000010001101000;
		weights[2508] <= 0000010111100011;
		weights[2509] <= 1000010001010111;
		weights[2510] <= 0000100010000011;
		weights[2511] <= 1000101101101100;
		weights[2512] <= 1001000110101110;
		weights[2513] <= 1000101010011110;
		weights[2514] <= 0000100001010110;
		weights[2515] <= 0000000001110110;
		weights[2516] <= 0000011000101001;
		weights[2517] <= 1000010011101010;
		weights[2518] <= 1000000000101010;
		weights[2519] <= 0000101011110011;
		weights[2520] <= 1000100011001110;
		weights[2521] <= 0000010010101100;
		weights[2522] <= 1000011010010111;
		weights[2523] <= 0000011101011110;
		weights[2524] <= 0000010101111100;
		weights[2525] <= 0000000110010010;
		weights[2526] <= 1000000001101001;
		weights[2527] <= 1000101110100100;
		weights[2528] <= 0000101001111101;
		weights[2529] <= 0000001001101000;
		weights[2530] <= 0000000010001100;
		weights[2531] <= 0000010011010000;
		weights[2532] <= 1000011110000001;
		weights[2533] <= 0000001011000101;
		weights[2534] <= 1000000000001010;
		weights[2535] <= 0000000100100000;
		weights[2536] <= 1000000110010110;
		weights[2537] <= 0000011110001001;
		weights[2538] <= 0000100011101010;
		weights[2539] <= 1000100000100101;
		weights[2540] <= 1000001111011001;
		weights[2541] <= 1000101110010001;
		weights[2542] <= 1000000100000010;
		weights[2543] <= 1000000010001001;
		weights[2544] <= 1000000101010001;
		weights[2545] <= 0000100001010010;
		weights[2546] <= 0000011110011101;
		weights[2547] <= 0000100010010110;
		weights[2548] <= 0000100000001001;
		weights[2549] <= 0001011000101001;
		weights[2550] <= 0000001111111110;
		weights[2551] <= 0000100001000101;
		weights[2552] <= 0000100011011010;
		weights[2553] <= 0000010000010001;
		weights[2554] <= 0000010111011011;
		weights[2555] <= 0000000101010011;
		weights[2556] <= 0000110001110000;
		weights[2557] <= 0000001110101011;
		weights[2558] <= 0000010001100110;
		weights[2559] <= 0000001010111010;
		weights[2560] <= 1000000011100011;
		weights[2561] <= 0000010101101101;
		weights[2562] <= 0000000111001110;
		weights[2563] <= 0000001100101111;
		weights[2564] <= 1000011001110111;
		weights[2565] <= 0000010111001001;
		weights[2566] <= 0000000100100010;
		weights[2567] <= 0000000011100001;
		weights[2568] <= 0000001110101011;
		weights[2569] <= 1000011110001011;
		weights[2570] <= 1000010110101011;
		weights[2571] <= 0000100001001000;
		weights[2572] <= 0000000000001000;
		weights[2573] <= 0000011101000111;
		weights[2574] <= 0000011000001110;
		weights[2575] <= 0000111001111011;
		weights[2576] <= 0000100000010101;
		weights[2577] <= 0000010001111011;
		weights[2578] <= 0001000110100001;
		weights[2579] <= 1000010101000111;
		weights[2580] <= 1000000001001100;
		weights[2581] <= 0000010100100010;
		weights[2582] <= 1001001000110000;
		weights[2583] <= 1000010111100110;
		weights[2584] <= 1000011010111001;
		weights[2585] <= 0000100100110011;
		weights[2586] <= 0000100101011010;
		weights[2587] <= 1000000100001000;
		weights[2588] <= 1000101011101101;
		weights[2589] <= 0000101111110110;
		weights[2590] <= 1000011000001000;
		weights[2591] <= 0001001001101000;
		weights[2592] <= 0000101011100111;
		weights[2593] <= 0000011001001110;
		weights[2594] <= 0000101100001010;
		weights[2595] <= 0000011010100000;
		weights[2596] <= 0000101000100110;
		weights[2597] <= 0000001011100010;
		weights[2598] <= 0000011100111101;
		weights[2599] <= 0001000011001011;
		weights[2600] <= 1000001110110010;
		weights[2601] <= 1000001100010110;
		weights[2602] <= 0000000000100001;
		weights[2603] <= 0000001010010110;
		weights[2604] <= 1000001010100111;
		weights[2605] <= 0000000010101111;
		weights[2606] <= 1000111001001001;
		weights[2607] <= 1000101011000011;
		weights[2608] <= 0000001010100001;
		weights[2609] <= 0000101100010111;
		weights[2610] <= 1000011101011111;
		weights[2611] <= 0000110011010011;
		weights[2612] <= 0000111110011100;
		weights[2613] <= 1000100111101010;
		weights[2614] <= 1000100111010010;
		weights[2615] <= 1000010111110100;
		weights[2616] <= 0000100100111101;
		weights[2617] <= 1000100101001100;
		weights[2618] <= 1000010011100010;
		weights[2619] <= 0000000110110101;
		weights[2620] <= 0000001000100010;
		weights[2621] <= 1000001110010101;
		weights[2622] <= 0000100011100100;
		weights[2623] <= 1000010011111100;
		weights[2624] <= 1000000001000011;
		weights[2625] <= 1000000101101010;
		weights[2626] <= 1000001111011111;
		weights[2627] <= 1000010100000110;
		weights[2628] <= 0000100001010100;
		weights[2629] <= 1000100110100000;
		weights[2630] <= 0000101010110111;
		weights[2631] <= 0000111000111011;
		weights[2632] <= 0000010001010110;
		weights[2633] <= 1000011100000010;
		weights[2634] <= 1000100010001111;
		weights[2635] <= 1000000011100000;
		weights[2636] <= 1000010101101010;
		weights[2637] <= 1001001000011111;
		weights[2638] <= 1000010101100111;
		weights[2639] <= 0000010011101010;
		weights[2640] <= 0000100100101101;
		weights[2641] <= 0000101110101110;
		weights[2642] <= 0000100100110011;
		weights[2643] <= 0000001010111000;
		weights[2644] <= 0000100111110110;
		weights[2645] <= 1000001111110010;
		weights[2646] <= 0000010011000000;
		weights[2647] <= 0000100011001001;
		weights[2648] <= 1000001001001110;
		weights[2649] <= 1000100100011110;
		weights[2650] <= 1001000101000111;
		weights[2651] <= 1000011100100101;
		weights[2652] <= 0000110001100100;
		weights[2653] <= 1000011001100000;
		weights[2654] <= 0000001000111110;
		weights[2655] <= 1000000010100111;
		weights[2656] <= 1000011101001111;
		weights[2657] <= 0000011000101010;
		weights[2658] <= 0000000000011001;
		weights[2659] <= 0000100010001101;
		weights[2660] <= 1000000010011010;
		weights[2661] <= 0000000011011110;
		weights[2662] <= 0000111010001001;
		weights[2663] <= 0000011101000010;
		weights[2664] <= 1000010111101101;
		weights[2665] <= 0000111111001101;
		weights[2666] <= 1000101000000100;
		weights[2667] <= 1000101010111010;
		weights[2668] <= 1000101101000011;
		weights[2669] <= 0000001011001000;
		weights[2670] <= 1000001001101101;
		weights[2671] <= 0000001101111010;
		weights[2672] <= 1000001010110010;
		weights[2673] <= 0000000110100101;
		weights[2674] <= 1000100010101001;
		weights[2675] <= 1000100110101111;
		weights[2676] <= 1000011111101111;
		weights[2677] <= 1000010111110100;
		weights[2678] <= 0000010110010000;
		weights[2679] <= 0000101011110001;
		weights[2680] <= 1000011110100000;
		weights[2681] <= 0000011101001101;
		weights[2682] <= 1000001110111101;
		weights[2683] <= 1000111111000111;
		weights[2684] <= 1000010101101111;
		weights[2685] <= 1000010101011010;
		weights[2686] <= 0000011010000101;
		weights[2687] <= 1000100100111010;
		weights[2688] <= 1000101000000011;
		weights[2689] <= 0000011001001010;
		weights[2690] <= 1001100000111101;
		weights[2691] <= 1000100001011000;
		weights[2692] <= 0000100110110100;
		weights[2693] <= 1000000010010000;
		weights[2694] <= 1000010010101110;
		weights[2695] <= 1000101110101001;
		weights[2696] <= 1000011101110110;
		weights[2697] <= 1000001101100011;
		weights[2698] <= 0001001010011101;
		weights[2699] <= 0000100101011101;
		weights[2700] <= 1000110100001011;
		weights[2701] <= 1000000000100100;
		weights[2702] <= 0000011000011001;
		weights[2703] <= 0000010111110011;
		weights[2704] <= 0000101000111000;
		weights[2705] <= 1000101011000010;
		weights[2706] <= 1000000001101000;
		weights[2707] <= 1000011011010010;
		weights[2708] <= 0000000110010000;
		weights[2709] <= 1000011000110101;
		weights[2710] <= 1000010101111000;
		weights[2711] <= 0000101000001001;
		weights[2712] <= 1000000110010010;
		weights[2713] <= 0000000111111000;
		weights[2714] <= 1000001111011100;
		weights[2715] <= 1000000100001011;
		weights[2716] <= 0000100000100111;
		weights[2717] <= 0000010011000100;
		weights[2718] <= 1000011100100101;
		weights[2719] <= 1000001101001011;
		weights[2720] <= 1000010010001001;
		weights[2721] <= 0000100000101100;
		weights[2722] <= 1000000010101001;
		weights[2723] <= 1000101110101100;
		weights[2724] <= 1001001010110110;
		weights[2725] <= 0000111001111000;
		weights[2726] <= 1000100101101100;
		weights[2727] <= 0000011001111101;
		weights[2728] <= 0000000010110001;
		weights[2729] <= 0000100001100110;
		weights[2730] <= 0001000000110011;
		weights[2731] <= 0000000110100000;
		weights[2732] <= 1000001111000011;
		weights[2733] <= 0000010001111011;
		weights[2734] <= 0000100001010100;
		weights[2735] <= 0000101111110100;
		weights[2736] <= 0000110001000000;
		weights[2737] <= 1000011001000111;
		weights[2738] <= 1000010110101010;
		weights[2739] <= 1000000001110010;
		weights[2740] <= 0000010100010000;
		weights[2741] <= 1000111001101100;
		weights[2742] <= 1000100000111000;
		weights[2743] <= 1000000100111101;
		weights[2744] <= 1000100100110000;
		weights[2745] <= 1000001110101101;
		weights[2746] <= 0000001011001100;
		weights[2747] <= 1000000011110010;
		weights[2748] <= 0000111101100011;
		weights[2749] <= 0000001100011111;
		weights[2750] <= 1000000110011001;
		weights[2751] <= 0000010010010100;
		weights[2752] <= 0000010101110111;
		weights[2753] <= 1000101110111001;
		weights[2754] <= 1000111100000010;
		weights[2755] <= 0000001110001100;
		weights[2756] <= 1000010101011000;
		weights[2757] <= 1000011011011010;
		weights[2758] <= 0000000110100111;
		weights[2759] <= 1000000100001101;
		weights[2760] <= 1000000110110000;
		weights[2761] <= 0000010010101111;
		weights[2762] <= 0000001000000011;
		weights[2763] <= 1000010000011010;
		weights[2764] <= 0000011010101011;
		weights[2765] <= 1000001010101100;
		weights[2766] <= 0000000010110001;
		weights[2767] <= 0000101010111000;
		weights[2768] <= 0000001111111110;
		weights[2769] <= 0000101010001001;
		weights[2770] <= 1000000001010000;
		weights[2771] <= 0000100100100000;
		weights[2772] <= 1000110010010001;
		weights[2773] <= 1000000000010000;
		weights[2774] <= 0000010100011101;
		weights[2775] <= 1000011001100001;
		weights[2776] <= 0000010101010111;
		weights[2777] <= 1000000011010001;
		weights[2778] <= 1000101001010001;
		weights[2779] <= 0000101110011111;
		weights[2780] <= 0001000011000001;
		weights[2781] <= 1001000110100000;
		weights[2782] <= 0000100010000101;
		weights[2783] <= 1000001101010000;
		weights[2784] <= 0000010100100010;
		weights[2785] <= 1000000011111001;
		weights[2786] <= 1001001011111101;
		weights[2787] <= 0000000101001111;
		weights[2788] <= 0000010001100101;
		weights[2789] <= 1000010110001000;
		weights[2790] <= 0000100111111100;
		weights[2791] <= 0000000111000111;
		weights[2792] <= 1000001110001100;
		weights[2793] <= 1000110101011011;
		weights[2794] <= 0000100100010100;
		weights[2795] <= 1000000101011111;
		weights[2796] <= 0000001101001110;
		weights[2797] <= 0000000110100110;
		weights[2798] <= 1000000010000001;
		weights[2799] <= 1000011111010000;
		weights[2800] <= 1001000010000010;
		weights[2801] <= 0000000111101011;
		weights[2802] <= 1000100111100010;
		weights[2803] <= 1000000011001011;
		weights[2804] <= 1000010010101100;
		weights[2805] <= 0000100000110100;
		weights[2806] <= 1001101110001001;
		weights[2807] <= 1000001101011001;
		weights[2808] <= 1000000110111100;
		weights[2809] <= 1000000000111000;
		weights[2810] <= 1001001000011100;
		weights[2811] <= 1000001001011001;
		weights[2812] <= 1000000010101101;
		weights[2813] <= 1000001001010111;
		weights[2814] <= 1000010001110110;
		weights[2815] <= 1000011001010111;
		weights[2816] <= 0000000110011100;
		weights[2817] <= 0000010000101101;
		weights[2818] <= 0000001001010100;
		weights[2819] <= 1000000100011100;
		weights[2820] <= 1000001100100101;
		weights[2821] <= 1000000001101010;
		weights[2822] <= 0000001011011010;
		weights[2823] <= 0000101010111011;
		weights[2824] <= 1000000110011000;
		weights[2825] <= 0000011101100110;
		weights[2826] <= 0000001010011100;
		weights[2827] <= 0000100110011100;
		weights[2828] <= 1000000111001100;
		weights[2829] <= 0000011101000011;
		weights[2830] <= 0000101100011110;
		weights[2831] <= 0000100000101011;
		weights[2832] <= 1000011010010010;
		weights[2833] <= 0000000110001001;
		weights[2834] <= 1000111010010001;
		weights[2835] <= 1000010011010111;
		weights[2836] <= 1000001010100110;
		weights[2837] <= 1000110011110010;
		weights[2838] <= 1000001000101011;
		weights[2839] <= 0000110110101110;
		weights[2840] <= 1000111010011100;
		weights[2841] <= 1000011000101000;
		weights[2842] <= 0000000001011010;
		weights[2843] <= 0000010011011010;
		weights[2844] <= 0000100000110100;
		weights[2845] <= 1000010010110110;
		weights[2846] <= 1001000010000111;
		weights[2847] <= 0000001000101100;
		weights[2848] <= 1000100010000110;
		weights[2849] <= 0000001000000110;
		weights[2850] <= 1000010001101111;
		weights[2851] <= 1000101101011011;
		weights[2852] <= 1000010011010101;
		weights[2853] <= 1000110001011110;
		weights[2854] <= 0000001100001101;
		weights[2855] <= 0000001110110011;
		weights[2856] <= 0000011000000001;
		weights[2857] <= 0000110101000001;
		weights[2858] <= 1000000111001101;
		weights[2859] <= 0000100101111001;
		weights[2860] <= 0000011110101011;
		weights[2861] <= 0000010000111111;
		weights[2862] <= 1000011101000000;
		weights[2863] <= 0000010111101000;
		weights[2864] <= 0000000110010101;
		weights[2865] <= 1000100110001111;
		weights[2866] <= 0000100000000110;
		weights[2867] <= 1000011001111001;
		weights[2868] <= 1000010111110010;
		weights[2869] <= 0000001010100001;
		weights[2870] <= 0000000011011011;
		weights[2871] <= 1000010000001111;
		weights[2872] <= 0000101011010101;
		weights[2873] <= 0000000111110110;
		weights[2874] <= 1000000010010101;
		weights[2875] <= 0000000101111101;
		weights[2876] <= 0000100110001010;
		weights[2877] <= 0000000010110001;
		weights[2878] <= 1000110110101100;
		weights[2879] <= 1000100001111010;
		weights[2880] <= 0000001011110110;
		weights[2881] <= 1000000100010110;
		weights[2882] <= 1000001101101100;
		weights[2883] <= 1000001110100101;
		weights[2884] <= 1000000001011000;
		weights[2885] <= 0000000011001100;
		weights[2886] <= 1000001010101011;
		weights[2887] <= 0000000001111001;
		weights[2888] <= 0000000011001111;
		weights[2889] <= 0000000010011110;
		weights[2890] <= 0000000011000100;
		weights[2891] <= 0000001000110000;
		weights[2892] <= 0000100010110100;
		weights[2893] <= 1000101011001110;
		weights[2894] <= 1000101011001100;
		weights[2895] <= 1000101100010100;
		weights[2896] <= 1000010011111110;
		weights[2897] <= 0000010100111101;
		weights[2898] <= 1000001101011000;
		weights[2899] <= 0000010010100011;
		weights[2900] <= 0000001110000111;
		weights[2901] <= 1000010010110100;
		weights[2902] <= 1000110010000101;
		weights[2903] <= 0000000000111101;
		weights[2904] <= 1000110111101010;
		weights[2905] <= 1000100000011111;
		weights[2906] <= 1000100011111101;
		weights[2907] <= 0000010000011010;
		weights[2908] <= 0000000011010110;
		weights[2909] <= 0000011111001001;
		weights[2910] <= 1000011011100100;
		weights[2911] <= 1000011000110100;
		weights[2912] <= 1000001000010111;
		weights[2913] <= 1000001011101001;
		weights[2914] <= 1000100001001010;
		weights[2915] <= 0000001011100110;
		weights[2916] <= 0000001010110111;
		weights[2917] <= 0000000111001100;
		weights[2918] <= 0000010010001111;
		weights[2919] <= 0000100101110100;
		weights[2920] <= 1000011000010011;
		weights[2921] <= 1000101111100100;
		weights[2922] <= 1000110111011101;
		weights[2923] <= 1000010011110001;
		weights[2924] <= 0000000101100111;
		weights[2925] <= 0000100110111001;
		weights[2926] <= 0000110101110101;
		weights[2927] <= 1000100011110011;
		weights[2928] <= 1000101110000011;
		weights[2929] <= 0000111100010100;
		weights[2930] <= 1000010010001010;
		weights[2931] <= 1000010001111001;
		weights[2932] <= 1001000110110001;
		weights[2933] <= 1000001011111110;
		weights[2934] <= 1000000100100001;
		weights[2935] <= 0000001011111100;
		weights[2936] <= 0000011000100110;
		weights[2937] <= 0000010100111001;
		weights[2938] <= 0000100110111001;
		weights[2939] <= 0000100110000011;
		weights[2940] <= 0000000110000011;
		weights[2941] <= 0001110111101101;
		weights[2942] <= 1000000111111001;
		weights[2943] <= 1000011001010010;
		weights[2944] <= 1000000001011001;
		weights[2945] <= 1000011110111111;
		weights[2946] <= 1000010100110011;
		weights[2947] <= 1000011110000110;
		weights[2948] <= 0000010001010011;
		weights[2949] <= 0000001000111101;
		weights[2950] <= 0000001101101111;
		weights[2951] <= 1000101110011101;
		weights[2952] <= 1000011111001011;
		weights[2953] <= 0000000111110100;
		weights[2954] <= 0000011110100011;
		weights[2955] <= 0000101000011101;
		weights[2956] <= 0000011000111100;
		weights[2957] <= 0000110000100001;
		weights[2958] <= 0001101001010001;
		weights[2959] <= 0001110101110001;
		weights[2960] <= 0001000101000010;
		weights[2961] <= 0000000001001111;
		weights[2962] <= 0000000101010010;
		weights[2963] <= 1000010000100001;
		weights[2964] <= 0000100101100011;
		weights[2965] <= 1000001111001101;
		weights[2966] <= 0000010101111011;
		weights[2967] <= 1000101000100001;
		weights[2968] <= 1000011010100001;
		weights[2969] <= 0000010110001010;
		weights[2970] <= 1000001111101111;
		weights[2971] <= 0000000100010011;
		weights[2972] <= 0000011111110100;
		weights[2973] <= 0000101111111000;
		weights[2974] <= 0000000111101100;
		weights[2975] <= 1000001101100000;
		weights[2976] <= 1000001100111101;
		weights[2977] <= 0000111001010110;
		weights[2978] <= 0000000110100000;
		weights[2979] <= 1000100000000010;
		weights[2980] <= 0000111101010101;
		weights[2981] <= 0000110101111011;
		weights[2982] <= 0000110011111000;
		weights[2983] <= 1000111100110000;
		weights[2984] <= 0000011111100001;
		weights[2985] <= 1000000111110001;
		weights[2986] <= 1000100110110010;
		weights[2987] <= 1000100101011100;
		weights[2988] <= 0000001011010011;
		weights[2989] <= 1000001111000000;
		weights[2990] <= 0000100111101110;
		weights[2991] <= 1000000100001000;
		weights[2992] <= 0000010100010000;
		weights[2993] <= 0000010001111000;
		weights[2994] <= 0000000100110111;
		weights[2995] <= 1000001111101110;
		weights[2996] <= 1000000100001011;
		weights[2997] <= 0000001111011010;
		weights[2998] <= 1000000111010100;
		weights[2999] <= 1001000000100101;
		weights[3000] <= 1000010000011001;
		weights[3001] <= 0000000101010011;
		weights[3002] <= 0000010100001111;
		weights[3003] <= 0000100010110100;
		weights[3004] <= 0000000010001101;
		weights[3005] <= 0000100011000000;
		weights[3006] <= 0000011101011011;
		weights[3007] <= 1000000011001100;
		weights[3008] <= 0000000111000001;
		weights[3009] <= 0000000010111001;
		weights[3010] <= 1000011100110011;
		weights[3011] <= 0000001101001100;
		weights[3012] <= 0000100010101100;
		weights[3013] <= 0000010001110001;
		weights[3014] <= 1000000011011010;
		weights[3015] <= 1000001101000100;
		weights[3016] <= 1000001001001011;
		weights[3017] <= 1000010110111011;
		weights[3018] <= 1000100001111000;
		weights[3019] <= 1000010110000000;
		weights[3020] <= 0000010100001101;
		weights[3021] <= 1000000100110000;
		weights[3022] <= 0000000101000000;
		weights[3023] <= 0000010001001001;
		weights[3024] <= 1000010001001010;
		weights[3025] <= 0000101000000010;
		weights[3026] <= 0000000011010111;
		weights[3027] <= 1000100011011110;
		weights[3028] <= 1000000100101010;
		weights[3029] <= 0000011000110010;
		weights[3030] <= 0000111000000100;
		weights[3031] <= 1000100101011001;
		weights[3032] <= 0000010010001001;
		weights[3033] <= 1000000001001000;
		weights[3034] <= 1000000101111001;
		weights[3035] <= 1000010101000001;
		weights[3036] <= 0000000000101011;
		weights[3037] <= 0000000000101111;
		weights[3038] <= 0000000000001001;
		weights[3039] <= 0000001010110011;
		weights[3040] <= 0000010101001110;
		weights[3041] <= 0000000001100011;
		weights[3042] <= 1000101011010100;
		weights[3043] <= 1000001010001010;
		weights[3044] <= 1000011000000001;
		weights[3045] <= 1000001010100110;
		weights[3046] <= 1000001100010001;
		weights[3047] <= 1000000100000111;
		weights[3048] <= 0000000110000111;
		weights[3049] <= 1000100000000101;
		weights[3050] <= 1000010111011110;
		weights[3051] <= 1000101111011001;
		weights[3052] <= 1000110110100100;
		weights[3053] <= 0000000010100110;
		weights[3054] <= 0000000001000000;
		weights[3055] <= 1000100010001001;
		weights[3056] <= 1000000000010010;
		weights[3057] <= 0000000010001111;
		weights[3058] <= 1000001000001000;
		weights[3059] <= 0000010001001101;
		weights[3060] <= 0000100001011110;
		weights[3061] <= 0000010101010110;
		weights[3062] <= 0000101010111000;
		weights[3063] <= 1000010111111111;
		weights[3064] <= 0000010110100001;
		weights[3065] <= 1000010110111100;
		weights[3066] <= 0000000001100110;
		weights[3067] <= 0000000000000100;
		weights[3068] <= 0000001100001000;
		weights[3069] <= 1000010100101101;
		weights[3070] <= 1000011001110101;
		weights[3071] <= 1000001010100000;
		weights[3072] <= 1000001011110100;
		weights[3073] <= 1000010000111001;
		weights[3074] <= 1000010000110111;
		weights[3075] <= 1000001000011100;
		weights[3076] <= 1000100111010110;
		weights[3077] <= 1000001100000001;
		weights[3078] <= 1000010011011100;
		weights[3079] <= 1000000011111100;
		weights[3080] <= 0000110001011100;
		weights[3081] <= 0000010101111100;
		weights[3082] <= 0000100010010101;
		weights[3083] <= 1000001100100111;
		weights[3084] <= 1000010000101101;
		weights[3085] <= 1000101001101101;
		weights[3086] <= 1000011110011110;
		weights[3087] <= 0000100100101010;
		weights[3088] <= 1000001110010000;
		weights[3089] <= 0000101111011010;
		weights[3090] <= 1000100000000101;
		weights[3091] <= 0000101111001100;
		weights[3092] <= 1000011000001011;
		weights[3093] <= 1000001011001111;
		weights[3094] <= 0000010111010000;
		weights[3095] <= 0000010001101100;
		weights[3096] <= 1000001011110001;
		weights[3097] <= 1000101111111011;
		weights[3098] <= 1000010000111011;
		weights[3099] <= 1000010000011111;
		weights[3100] <= 1000010001001001;
		weights[3101] <= 1000001010101101;
		weights[3102] <= 0000101010011011;
		weights[3103] <= 0000010000000110;
		weights[3104] <= 1000001000110011;
		weights[3105] <= 1000110001101110;
		weights[3106] <= 0000000110001011;
		weights[3107] <= 1000011000000111;
		weights[3108] <= 0000001001111000;
		weights[3109] <= 1000001010000000;
		weights[3110] <= 0001010010010010;
		weights[3111] <= 1000110011011101;
		weights[3112] <= 0000011101000011;
		weights[3113] <= 0000001110001101;
		weights[3114] <= 1000010111100010;
		weights[3115] <= 0000110011101110;
		weights[3116] <= 1000010111000100;
		weights[3117] <= 1000010110010001;
		weights[3118] <= 1001000101011110;
		weights[3119] <= 0000011110100110;
		weights[3120] <= 0000001100000001;
		weights[3121] <= 1000100000101001;
		weights[3122] <= 0000011001000001;
		weights[3123] <= 1000000111011101;
		weights[3124] <= 1001010000001011;
		weights[3125] <= 0000011001110100;
		weights[3126] <= 1000110010101111;
		weights[3127] <= 1000011111001000;
		weights[3128] <= 1000001101111110;
		weights[3129] <= 0000001111010100;
		weights[3130] <= 0000010100110001;
		weights[3131] <= 0000000000111000;
		weights[3132] <= 0000011110000010;
		weights[3133] <= 0000101000110001;
		weights[3134] <= 1000010001000111;
		weights[3135] <= 1000000000101000;
		weights[3136] <= 1000000011000010;
		weights[3137] <= 1000001100001110;
		weights[3138] <= 1000011011110111;
		weights[3139] <= 1000100010101001;
		weights[3140] <= 0001000110001010;
		weights[3141] <= 1000000010110101;
		weights[3142] <= 0000101101111010;
		weights[3143] <= 1000000000110001;
		weights[3144] <= 0000101001000111;
		weights[3145] <= 1000001110110001;
		weights[3146] <= 1001001100111001;
		weights[3147] <= 0000101110110001;
		weights[3148] <= 1000000010110100;
		weights[3149] <= 0001010010111110;
		weights[3150] <= 1000000110111001;
		weights[3151] <= 1000010100101011;
		weights[3152] <= 0000100001011000;
		weights[3153] <= 1000100010110011;
		weights[3154] <= 1000110111110101;
		weights[3155] <= 0000010101010101;
		weights[3156] <= 0000011010101011;
		weights[3157] <= 1000100110000101;
		weights[3158] <= 0000010110110111;
		weights[3159] <= 1000001101111011;
		weights[3160] <= 0001000100000010;
		weights[3161] <= 0000000111101110;
		weights[3162] <= 0000111001100001;
		weights[3163] <= 0001001100110111;
		weights[3164] <= 0000010111001100;
		weights[3165] <= 1000100000100111;
		weights[3166] <= 1000110001100011;
		weights[3167] <= 1000010110000001;
		weights[3168] <= 1000000011101110;
		weights[3169] <= 1000011010011011;
		weights[3170] <= 1000111010010001;
		weights[3171] <= 0000100101101101;
		weights[3172] <= 0000010000001100;
		weights[3173] <= 0000000011000101;
		weights[3174] <= 0001010000011100;
		weights[3175] <= 1000001010011000;
		weights[3176] <= 1000110000100000;
		weights[3177] <= 0000100000100110;
		weights[3178] <= 1000001101101110;
		weights[3179] <= 0000110000101101;
		weights[3180] <= 1000100000111111;
		weights[3181] <= 0000001010000110;
		weights[3182] <= 1001100100101000;
		weights[3183] <= 1000011011000111;
		weights[3184] <= 1000010011101100;
		weights[3185] <= 0000010100100100;
		weights[3186] <= 1001000111101111;
		weights[3187] <= 1000001100000101;
		weights[3188] <= 0000100101111111;
		weights[3189] <= 0001000000000010;
		weights[3190] <= 1000011001100011;
		weights[3191] <= 0000001010010001;
		weights[3192] <= 0000101011100110;
		weights[3193] <= 1000010101101101;
		weights[3194] <= 0000011011100110;
		weights[3195] <= 1000001100101101;
		weights[3196] <= 1000010000011001;
		weights[3197] <= 1000001010100101;
		weights[3198] <= 1000010111011001;
		weights[3199] <= 0000110011111110;
		weights[3200] <= 1000110000011001;
		weights[3201] <= 1000001011111001;
		weights[3202] <= 0000010000011111;
		weights[3203] <= 1000100110011010;
		weights[3204] <= 0000000100000000;
		weights[3205] <= 1000001100111100;
		weights[3206] <= 1000010001101111;
		weights[3207] <= 0000001001011100;
		weights[3208] <= 1000000100101001;
		weights[3209] <= 0000011100010110;
		weights[3210] <= 0000011001001111;
		weights[3211] <= 1000001011100100;
		weights[3212] <= 0000000001100101;
		weights[3213] <= 0000011100001101;
		weights[3214] <= 0000000010010001;
		weights[3215] <= 0000001110110001;
		weights[3216] <= 0000100011111001;
		weights[3217] <= 1000000111010001;
		weights[3218] <= 1000101110111101;
		weights[3219] <= 1000001010011000;
		weights[3220] <= 1000100101111010;
		weights[3221] <= 1000001111001111;
		weights[3222] <= 1000001010010111;
		weights[3223] <= 0000000100100111;
		weights[3224] <= 0000100000100110;
		weights[3225] <= 0000011001010001;
		weights[3226] <= 0000000001111100;
		weights[3227] <= 1000000100000001;
		weights[3228] <= 1000001110010001;
		weights[3229] <= 1000001010001011;
		weights[3230] <= 1000011001001101;
		weights[3231] <= 0000000011111101;
		weights[3232] <= 1000101111101001;
		weights[3233] <= 1000111001110110;
		weights[3234] <= 0000010011110000;
		weights[3235] <= 0000100011110111;
		weights[3236] <= 0000010010010001;
		weights[3237] <= 0000111110000111;
		weights[3238] <= 1000111110010111;
		weights[3239] <= 1000001011011111;
		weights[3240] <= 1000000000010001;
		weights[3241] <= 0000010111001100;
		weights[3242] <= 0000101000100100;
		weights[3243] <= 1000011110010010;
		weights[3244] <= 1000100110000001;
		weights[3245] <= 0000101000100111;
		weights[3246] <= 1000001001010110;
		weights[3247] <= 0000001000001111;
		weights[3248] <= 0000000101000000;
		weights[3249] <= 1000110010010100;
		weights[3250] <= 1000001110101001;
		weights[3251] <= 0000011000110001;
		weights[3252] <= 1000100110010011;
		weights[3253] <= 1000100110001001;
		weights[3254] <= 1000011011010000;
		weights[3255] <= 0000101110111101;
		weights[3256] <= 0000110111011100;
		weights[3257] <= 1000000110011100;
		weights[3258] <= 1000000000001101;
		weights[3259] <= 1000101001111101;
		weights[3260] <= 0000000110101010;
		weights[3261] <= 0000010011110000;
		weights[3262] <= 1000000001010010;
		weights[3263] <= 0000001000100011;
		weights[3264] <= 1000110011100111;
		weights[3265] <= 1000011101010101;
		weights[3266] <= 1000010111100011;
		weights[3267] <= 1000000000110111;
		weights[3268] <= 1000011100000110;
		weights[3269] <= 1000000111010000;
		weights[3270] <= 1000010001100010;
		weights[3271] <= 0000010111011110;
		weights[3272] <= 0000000000110011;
		weights[3273] <= 0001010011000110;
		weights[3274] <= 0000100111111101;
		weights[3275] <= 1000001000110111;
		weights[3276] <= 1000011101011000;
		weights[3277] <= 0000011011111000;
		weights[3278] <= 1000100011101010;
		weights[3279] <= 1000110100011010;
		weights[3280] <= 1000000101011111;
		weights[3281] <= 0000001111101100;
		weights[3282] <= 0000001000110001;
		weights[3283] <= 0000001110010001;
		weights[3284] <= 1000000110101011;
		weights[3285] <= 0000001111000010;
		weights[3286] <= 1000100000111001;
		weights[3287] <= 0000001101001011;
		weights[3288] <= 0000000000000101;
		weights[3289] <= 1000000000011000;
		weights[3290] <= 1000100000010100;
		weights[3291] <= 0000101010010011;
		weights[3292] <= 0000010111100000;
		weights[3293] <= 0001001001110110;
		weights[3294] <= 0000101111110011;
		weights[3295] <= 0000001010101100;
		weights[3296] <= 1000001011001101;
		weights[3297] <= 0000011011011010;
		weights[3298] <= 0000010111100111;
		weights[3299] <= 1000100010100101;
		weights[3300] <= 1000001010001001;
		weights[3301] <= 1000100011110100;
		weights[3302] <= 0000010011110100;
		weights[3303] <= 1000100111010011;
		weights[3304] <= 1000010100010100;
		weights[3305] <= 0000111110001100;
		weights[3306] <= 1000100100111000;
		weights[3307] <= 1000100011111001;
		weights[3308] <= 1000010001110011;
		weights[3309] <= 1000111000010010;
		weights[3310] <= 1000011101100001;
		weights[3311] <= 1000101101001000;
		weights[3312] <= 1000100011101100;
		weights[3313] <= 0000000001001101;
		weights[3314] <= 0000000101110110;
		weights[3315] <= 1000111000011000;
		weights[3316] <= 0000100000101111;
		weights[3317] <= 0000010001101101;
		weights[3318] <= 0000001110000000;
		weights[3319] <= 0000000001110110;
		weights[3320] <= 0000101010110010;
		weights[3321] <= 0000010100110100;
		weights[3322] <= 0000001001110110;
		weights[3323] <= 1000110000100010;
		weights[3324] <= 0000011000100101;
		weights[3325] <= 0000101000010111;
		weights[3326] <= 0000000000010100;
		weights[3327] <= 1000000100101000;
		weights[3328] <= 0000000111100110;
		weights[3329] <= 0000001111000011;
		weights[3330] <= 0000000110111011;
		weights[3331] <= 0000000110001110;
		weights[3332] <= 1000010100110101;
		weights[3333] <= 1000011111110000;
		weights[3334] <= 1000101000100110;
		weights[3335] <= 1000111100100100;
		weights[3336] <= 1000100101000001;
		weights[3337] <= 1000000111011001;
		weights[3338] <= 0000001001010001;
		weights[3339] <= 1000000010100100;
		weights[3340] <= 0000100000101111;
		weights[3341] <= 0000111100101010;
		weights[3342] <= 0000101011011000;
		weights[3343] <= 1000111011010001;
		weights[3344] <= 1001000010100001;
		weights[3345] <= 1000110001000111;
		weights[3346] <= 1000011110001100;
		weights[3347] <= 0000011111001101;
		weights[3348] <= 0000100110110001;
		weights[3349] <= 0000001010111100;
		weights[3350] <= 0000011011110010;
		weights[3351] <= 0000011000101001;
		weights[3352] <= 0000100110010000;
		weights[3353] <= 1000010010101010;
		weights[3354] <= 1000010101111111;
		weights[3355] <= 1000110111010110;
		weights[3356] <= 1000011000110000;
		weights[3357] <= 1000100110100101;
		weights[3358] <= 0000001010101100;
		weights[3359] <= 0000010110110001;
		weights[3360] <= 0000110100111010;
		weights[3361] <= 0000000101010011;
		weights[3362] <= 0001101101000000;
		weights[3363] <= 0000111011010011;
		weights[3364] <= 1000000001100100;
		weights[3365] <= 1000000010111001;
		weights[3366] <= 0000110101100100;
		weights[3367] <= 1000100010100001;
		weights[3368] <= 0000010011110101;
		weights[3369] <= 0000000110111111;
		weights[3370] <= 0001010001001110;
		weights[3371] <= 1000001000011111;
		weights[3372] <= 0000001001101000;
		weights[3373] <= 0000011011010111;
		weights[3374] <= 1000010001100001;
		weights[3375] <= 1000011100100100;
		weights[3376] <= 1000000010011111;
		weights[3377] <= 0000100001110000;
		weights[3378] <= 0000010010100001;
		weights[3379] <= 1000001110101100;
		weights[3380] <= 0000100101010011;
		weights[3381] <= 0000110011101100;
		weights[3382] <= 0000011001100110;
		weights[3383] <= 1000000110110111;
		weights[3384] <= 0000011111011000;
		weights[3385] <= 0000100010101110;
		weights[3386] <= 1000011110010111;
		weights[3387] <= 0000100011000110;
		weights[3388] <= 1000010110110100;
		weights[3389] <= 1000011110010110;
		weights[3390] <= 1000001010100001;
		weights[3391] <= 0000011101000001;
		weights[3392] <= 1001001011011101;
		weights[3393] <= 0000001000100100;
		weights[3394] <= 0000011110100101;
		weights[3395] <= 1000000010011101;
		weights[3396] <= 0001010100110001;
		weights[3397] <= 0000010110101100;
		weights[3398] <= 0000101000100000;
		weights[3399] <= 1000010111001011;
		weights[3400] <= 1000101011000101;
		weights[3401] <= 1000001011010101;
		weights[3402] <= 1000001011100100;
		weights[3403] <= 1000000011010001;
		weights[3404] <= 0000011110010111;
		weights[3405] <= 0000001110011010;
		weights[3406] <= 0000100011101011;
		weights[3407] <= 0000100000101001;
		weights[3408] <= 1000010010110000;
		weights[3409] <= 0000000100001110;
		weights[3410] <= 0000011011010110;
		weights[3411] <= 0000110100101100;
		weights[3412] <= 0000000110001111;
		weights[3413] <= 1000001100001011;
		weights[3414] <= 0000010101100100;
		weights[3415] <= 0000100111110111;
		weights[3416] <= 1000001101010000;
		weights[3417] <= 1000100100100110;
		weights[3418] <= 1001000100101011;
		weights[3419] <= 1000110110010110;
		weights[3420] <= 1000100011101111;
		weights[3421] <= 1000001001110110;
		weights[3422] <= 1000000101100111;
		weights[3423] <= 1000111000011111;
		weights[3424] <= 1000111110010100;
		weights[3425] <= 1000010101111001;
		weights[3426] <= 1000101101010100;
		weights[3427] <= 0000010101001001;
		weights[3428] <= 0000001011101000;
		weights[3429] <= 1000010001001100;
		weights[3430] <= 1000011011101101;
		weights[3431] <= 1000010011000101;
		weights[3432] <= 0000000000110101;
		weights[3433] <= 1000011000000101;
		weights[3434] <= 1000000011011110;
		weights[3435] <= 0000100101111011;
		weights[3436] <= 0000010100110111;
		weights[3437] <= 1000101111010100;
		weights[3438] <= 1000110110001101;
		weights[3439] <= 1000001100010011;
		weights[3440] <= 0000000100001000;
		weights[3441] <= 1000010111101000;
		weights[3442] <= 1000000111010000;
		weights[3443] <= 1000001111000001;
		weights[3444] <= 1000000011100100;
		weights[3445] <= 1000110111100010;
		weights[3446] <= 0000001000110100;
		weights[3447] <= 1000010101000011;
		weights[3448] <= 1000010011010001;
		weights[3449] <= 0000100010111011;
		weights[3450] <= 1000000001000010;
		weights[3451] <= 1000000011111011;
		weights[3452] <= 1000011100001011;
		weights[3453] <= 1000011000101100;
		weights[3454] <= 1000001101001010;
		weights[3455] <= 0000000100100001;
		weights[3456] <= 0000111111001001;
		weights[3457] <= 0000000100110001;
		weights[3458] <= 0000010100000001;
		weights[3459] <= 0000110101011111;
		weights[3460] <= 1000001111110100;
		weights[3461] <= 0000000010101000;
		weights[3462] <= 1000001101001011;
		weights[3463] <= 1000000010111100;
		weights[3464] <= 1000001000110110;
		weights[3465] <= 0000011010001001;
		weights[3466] <= 0000001110010001;
		weights[3467] <= 0000000101101011;
		weights[3468] <= 1001000011100100;
		weights[3469] <= 1000010001101000;
		weights[3470] <= 0000100000110100;
		weights[3471] <= 0000001101000110;
		weights[3472] <= 1000101111101011;
		weights[3473] <= 1000001000101100;
		weights[3474] <= 0000000011000100;
		weights[3475] <= 0000000110001101;
		weights[3476] <= 0000101011000101;
		weights[3477] <= 0000110111111111;
		weights[3478] <= 0000100101110101;
		weights[3479] <= 1000001110001101;
		weights[3480] <= 0000000010000111;
		weights[3481] <= 0000001101100111;
		weights[3482] <= 1000011000001111;
		weights[3483] <= 0000000111001111;
		weights[3484] <= 0000011111100010;
		weights[3485] <= 1000011101011001;
		weights[3486] <= 0000101011101110;
		weights[3487] <= 0000010001101011;
		weights[3488] <= 0000001111010001;
		weights[3489] <= 0000101001101010;
		weights[3490] <= 1000010011010000;
		weights[3491] <= 0000000111111010;
		weights[3492] <= 1000010111111010;
		weights[3493] <= 0000110000001100;
		weights[3494] <= 0000001010111111;
		weights[3495] <= 1000010011010110;
		weights[3496] <= 1000010011111101;
		weights[3497] <= 0000001111101011;
		weights[3498] <= 1000000111011111;
		weights[3499] <= 1000010011001100;
		weights[3500] <= 0000011100111101;
		weights[3501] <= 1000001000110011;
		weights[3502] <= 1000010010000100;
		weights[3503] <= 0000101100000000;
		weights[3504] <= 1000001111101001;
		weights[3505] <= 1000001101011000;
		weights[3506] <= 1000001001100010;
		weights[3507] <= 0000100110000000;
		weights[3508] <= 1000010011000111;
		weights[3509] <= 0000110100010011;
		weights[3510] <= 0000100011001100;
		weights[3511] <= 0000001111100111;
		weights[3512] <= 1000111011001000;
		weights[3513] <= 1000110010101110;
		weights[3514] <= 0000011011000100;
		weights[3515] <= 0000000100101011;
		weights[3516] <= 0000011101110100;
		weights[3517] <= 1000011010110111;
		weights[3518] <= 1000100101001011;
		weights[3519] <= 0000011100001111;
		weights[3520] <= 0000010111001000;
		weights[3521] <= 1000010011011100;
		weights[3522] <= 1000110000101000;
		weights[3523] <= 0000001110001101;
		weights[3524] <= 1000000111011010;
		weights[3525] <= 1000001100111110;
		weights[3526] <= 1000011001010000;
		weights[3527] <= 0000100111101010;
		weights[3528] <= 0000100110110100;
		weights[3529] <= 0000011001001100;
		weights[3530] <= 1000100100100011;
		weights[3531] <= 1000100111101110;
		weights[3532] <= 1000001000100000;
		weights[3533] <= 1001010000100111;
		weights[3534] <= 0000000001011100;
		weights[3535] <= 0000000111011000;
		weights[3536] <= 0000010000000000;
		weights[3537] <= 0000001010000001;
		weights[3538] <= 0000010001011011;
		weights[3539] <= 0000010111100001;
		weights[3540] <= 0000111000001000;
		weights[3541] <= 0000001111110110;
		weights[3542] <= 1000101111110011;
		weights[3543] <= 1000011111100100;
		weights[3544] <= 0000110010111001;
		weights[3545] <= 1000010010111011;
		weights[3546] <= 0000000011000111;
		weights[3547] <= 0000010001001111;
		weights[3548] <= 0000100011111001;
		weights[3549] <= 1000010100110101;
		weights[3550] <= 1000001011000110;
		weights[3551] <= 0000000101101010;
		weights[3552] <= 1000101011100111;
		weights[3553] <= 0000111001001111;
		weights[3554] <= 0000001100000000;
		weights[3555] <= 0000001000001100;
		weights[3556] <= 0000110101100001;
		weights[3557] <= 0001010011010000;
		weights[3558] <= 1000011011011011;
		weights[3559] <= 1000001100101111;
		weights[3560] <= 1000011110101110;
		weights[3561] <= 0000011011011001;
		weights[3562] <= 0000000100110100;
		weights[3563] <= 0000000101000110;
		weights[3564] <= 1000101001001001;
		weights[3565] <= 1000010010101000;
		weights[3566] <= 1000101000111000;
		weights[3567] <= 0000001001010111;
		weights[3568] <= 0000010100111010;
		weights[3569] <= 0000110010000001;
		weights[3570] <= 1000001110110001;
		weights[3571] <= 1000101010111100;
		weights[3572] <= 1000111000010110;
		weights[3573] <= 1001010100001010;
		weights[3574] <= 1000001010000011;
		weights[3575] <= 1000101101000100;
		weights[3576] <= 1000111110110010;
		weights[3577] <= 0000011100101101;
		weights[3578] <= 1000010001010100;
		weights[3579] <= 1000000101100010;
		weights[3580] <= 1000011010000011;
		weights[3581] <= 0000101111111110;
		weights[3582] <= 1000110011111010;
		weights[3583] <= 0000010000110011;
		weights[3584] <= 1000010000101010;
		weights[3585] <= 0000111001100000;
		weights[3586] <= 1000110100110101;
		weights[3587] <= 0000011110100000;
		weights[3588] <= 1000110100100001;
		weights[3589] <= 0000001100011111;
		weights[3590] <= 1000000000110100;
		weights[3591] <= 0000110011101010;
		weights[3592] <= 0000001000101010;
		weights[3593] <= 0000000110101000;
		weights[3594] <= 0000000001110001;
		weights[3595] <= 1000010001111100;
		weights[3596] <= 0000010010111011;
		weights[3597] <= 0000001001111101;
		weights[3598] <= 0000001110010000;
		weights[3599] <= 1000000010100111;
		weights[3600] <= 1001000001110001;
		weights[3601] <= 1000001001011111;
		weights[3602] <= 1000100010000011;
		weights[3603] <= 0000011010011001;
		weights[3604] <= 1000111001111011;
		weights[3605] <= 1000010100000001;
		weights[3606] <= 0000011100101011;
		weights[3607] <= 0000110110100100;
		weights[3608] <= 0000000011001111;
		weights[3609] <= 1000011010000111;
		weights[3610] <= 0000000010100010;
		weights[3611] <= 0000000110110110;
		weights[3612] <= 1000110100001001;
		weights[3613] <= 0000010101010101;
		weights[3614] <= 1000011110100110;
		weights[3615] <= 0000011000000110;
		weights[3616] <= 1000010100001110;
		weights[3617] <= 1000010111000110;
		weights[3618] <= 1000100110101111;
		weights[3619] <= 0000000101001000;
		weights[3620] <= 0000001011110101;
		weights[3621] <= 1000101011101111;
		weights[3622] <= 1000000110111010;
		weights[3623] <= 0000100010101101;
		weights[3624] <= 1000010011001100;
		weights[3625] <= 1000000010011010;
		weights[3626] <= 1000100011110010;
		weights[3627] <= 1000000000000001;
		weights[3628] <= 0000010111011010;
		weights[3629] <= 0000001000100010;
		weights[3630] <= 1000100000100100;
		weights[3631] <= 1001000101100011;
		weights[3632] <= 0000001110100100;
		weights[3633] <= 1000000111011011;
		weights[3634] <= 0000010111110000;
		weights[3635] <= 0000000011110111;
		weights[3636] <= 0001000101111011;
		weights[3637] <= 0000010000100000;
		weights[3638] <= 0000000010010110;
		weights[3639] <= 0000010100000111;
		weights[3640] <= 1000001010101010;
		weights[3641] <= 0000111100001111;
		weights[3642] <= 1000111001110110;
		weights[3643] <= 0000111101010111;
		weights[3644] <= 0000000010110011;
		weights[3645] <= 0000001010000000;
		weights[3646] <= 0001000110100110;
		weights[3647] <= 0000000101100011;
		weights[3648] <= 0001000001101011;
		weights[3649] <= 0000000110101010;
		weights[3650] <= 0000010101111100;
		weights[3651] <= 0000010111100010;
		weights[3652] <= 0000001110000000;
		weights[3653] <= 1000001001101000;
		weights[3654] <= 0000101001101110;
		weights[3655] <= 0000000111110001;
		weights[3656] <= 0000011110001011;
		weights[3657] <= 0000000000100011;
		weights[3658] <= 1000110001111000;
		weights[3659] <= 1000101101110100;
		weights[3660] <= 0000001101100001;
		weights[3661] <= 0000001010111111;
		weights[3662] <= 1000110111011110;
		weights[3663] <= 1000011010111101;
		weights[3664] <= 0000000011101111;
		weights[3665] <= 0000001111011100;
		weights[3666] <= 1000101000000011;
		weights[3667] <= 0000011001110001;
		weights[3668] <= 0000000100110000;
		weights[3669] <= 0000001010011000;
		weights[3670] <= 0000001011000001;
		weights[3671] <= 0000000101100100;
		weights[3672] <= 1000100100010110;
		weights[3673] <= 0000111110001101;
		weights[3674] <= 1000011000001100;
		weights[3675] <= 1000010110001011;
		weights[3676] <= 0000011101110110;
		weights[3677] <= 1000011001100101;
		weights[3678] <= 1000010101101010;
		weights[3679] <= 1000110000010111;
		weights[3680] <= 0000100100001010;
		weights[3681] <= 0000000010111110;
		weights[3682] <= 1000010001110010;
		weights[3683] <= 0000001011110100;
		weights[3684] <= 0000000100110110;
		weights[3685] <= 0000010001011001;
		weights[3686] <= 1000001000000001;
		weights[3687] <= 0000000001001001;
		weights[3688] <= 0000101011111110;
		weights[3689] <= 0000110111111011;
		weights[3690] <= 1000011111010010;
		weights[3691] <= 1000101100011011;
		weights[3692] <= 0000000000110100;
		weights[3693] <= 0000100110110011;
		weights[3694] <= 1000001100111110;
		weights[3695] <= 0000011110000001;
		weights[3696] <= 0000011000000010;
		weights[3697] <= 0000000110011001;
		weights[3698] <= 0000101011100000;
		weights[3699] <= 0000001110000011;
		weights[3700] <= 1000011001111110;
		weights[3701] <= 0000011101110100;
		weights[3702] <= 0000011100000011;
		weights[3703] <= 1000111111010110;
		weights[3704] <= 1000000010100110;
		weights[3705] <= 0000010000011110;
		weights[3706] <= 1000011110001111;
		weights[3707] <= 1000011010001100;
		weights[3708] <= 1000110010111110;
		weights[3709] <= 0000100000001000;
		weights[3710] <= 0000010101100001;
		weights[3711] <= 1000101110101101;
		weights[3712] <= 0000000011110110;
		weights[3713] <= 1000100110100010;
		weights[3714] <= 1000101100001000;
		weights[3715] <= 1000100100001101;
		weights[3716] <= 1000110011001001;
		weights[3717] <= 1000000001101100;
		weights[3718] <= 1000010100101011;
		weights[3719] <= 1000001100100011;
		weights[3720] <= 0000011100010011;
		weights[3721] <= 1000000010101011;
		weights[3722] <= 1000001010111010;
		weights[3723] <= 1000011110100010;
		weights[3724] <= 1000110011000110;
		weights[3725] <= 1001000101101100;
		weights[3726] <= 0000010111101011;
		weights[3727] <= 1000010111110001;
		weights[3728] <= 1000011110110001;
		weights[3729] <= 1000100011101111;
		weights[3730] <= 0000011111011001;
		weights[3731] <= 1000010110010111;
		weights[3732] <= 1000010001011111;
		weights[3733] <= 1000010111001100;
		weights[3734] <= 1000100001001110;
		weights[3735] <= 1000001100111011;
		weights[3736] <= 1000001010110110;
		weights[3737] <= 1000010100100111;
		weights[3738] <= 1000010100100011;
		weights[3739] <= 1000001000111110;
		weights[3740] <= 1000100000011100;
		weights[3741] <= 0000000010000011;
		weights[3742] <= 1000011111101110;
		weights[3743] <= 1000001110000010;
		weights[3744] <= 0000010011110100;
		weights[3745] <= 0000010100011101;
		weights[3746] <= 1000011010101100;
		weights[3747] <= 0000010000111000;
		weights[3748] <= 1000110011101000;
		weights[3749] <= 0000101110000101;
		weights[3750] <= 1000101001010001;
		weights[3751] <= 0000010011000111;
		weights[3752] <= 0000100110111001;
		weights[3753] <= 1000101010010011;
		weights[3754] <= 1000001000011101;
		weights[3755] <= 1000110100001000;
		weights[3756] <= 1000010101011101;
		weights[3757] <= 1000100000110011;
		weights[3758] <= 0000000110101000;
		weights[3759] <= 0000110010101100;
		weights[3760] <= 0000100101101100;
		weights[3761] <= 0000010100000011;
		weights[3762] <= 1000011000110111;
		weights[3763] <= 0000010010111111;
		weights[3764] <= 0000000111000101;
		weights[3765] <= 0000000111110011;
		weights[3766] <= 0000111000000010;
		weights[3767] <= 0000111010100010;
		weights[3768] <= 0000010000001111;
		weights[3769] <= 1000000101010001;
		weights[3770] <= 1000000011010111;
		weights[3771] <= 0000001000110100;
		weights[3772] <= 1001000011101011;
		weights[3773] <= 1000011000000111;
		weights[3774] <= 1000100111101010;
		weights[3775] <= 1000000110010010;
		weights[3776] <= 1001010101001000;
		weights[3777] <= 0000010000111100;
		weights[3778] <= 0001000101110001;
		weights[3779] <= 1000001010101010;
		weights[3780] <= 0000010111100100;
		weights[3781] <= 1000010101001111;
		weights[3782] <= 1000010101111011;
		weights[3783] <= 1000000111011001;
		weights[3784] <= 0000101011001001;
		weights[3785] <= 1000100001010101;
		weights[3786] <= 0000011001010000;
		weights[3787] <= 1000000100101100;
		weights[3788] <= 1000100110011000;
		weights[3789] <= 0000111100010111;
		weights[3790] <= 0000000010110101;
		weights[3791] <= 1000100110110100;
		weights[3792] <= 1000110110101000;
		weights[3793] <= 1000001111111111;
		weights[3794] <= 1000011101001101;
		weights[3795] <= 1000010101111110;
		weights[3796] <= 1000100000000101;
		weights[3797] <= 1000001110111010;
		weights[3798] <= 0000001101011100;
		weights[3799] <= 0000010111100101;
		weights[3800] <= 0000011110011001;
		weights[3801] <= 0000100010100110;
		weights[3802] <= 1000010111110010;
		weights[3803] <= 1000001011000011;
		weights[3804] <= 0000010000000000;
		weights[3805] <= 1000010000011011;
		weights[3806] <= 1000001000011011;
		weights[3807] <= 0000100101010100;
		weights[3808] <= 1000000101011111;
		weights[3809] <= 0000101010100110;
		weights[3810] <= 0000000111010111;
		weights[3811] <= 1000000110011100;
		weights[3812] <= 1000100010111011;
		weights[3813] <= 0000101000111110;
		weights[3814] <= 0000001000010001;
		weights[3815] <= 0000000000000011;
		weights[3816] <= 1000010111101011;
		weights[3817] <= 0000010010101000;
		weights[3818] <= 0001001010010001;
		weights[3819] <= 0001000101101011;
		weights[3820] <= 0001010110001000;
		weights[3821] <= 0000100100001111;
		weights[3822] <= 1000001111100111;
		weights[3823] <= 0000010011011001;
		weights[3824] <= 0000000000110100;
		weights[3825] <= 0000101101111010;
		weights[3826] <= 1000000111110100;
		weights[3827] <= 1000010111110101;
		weights[3828] <= 0000000001010000;
		weights[3829] <= 0000101001011111;
		weights[3830] <= 0000001001101100;
		weights[3831] <= 0000100111010000;
		weights[3832] <= 0000001101101101;
		weights[3833] <= 0000011010000011;
		weights[3834] <= 0000011110100101;
		weights[3835] <= 0000010000101101;
		weights[3836] <= 1000101110111101;
		weights[3837] <= 1000010010011010;
		weights[3838] <= 0000110001011101;
		weights[3839] <= 0000110111100010;
		weights[3840] <= 0000010010100000;
		weights[3841] <= 1000001010011100;
		weights[3842] <= 0000011010101111;
		weights[3843] <= 0000001111111000;
		weights[3844] <= 1000011011000100;
		weights[3845] <= 0000000101100110;
		weights[3846] <= 1000100001111011;
		weights[3847] <= 0000010100101001;
		weights[3848] <= 0000101010111111;
		weights[3849] <= 1000010111000100;
		weights[3850] <= 0000000101100101;
		weights[3851] <= 0000010011010001;
		weights[3852] <= 1001000001100111;
		weights[3853] <= 0000100001110110;
		weights[3854] <= 0000000111110011;
		weights[3855] <= 0000011010100001;
		weights[3856] <= 1000101100000111;
		weights[3857] <= 1000011101010001;
		weights[3858] <= 1000010011010101;
		weights[3859] <= 0000011101111111;
		weights[3860] <= 1000000101100101;
		weights[3861] <= 0000011011111110;
		weights[3862] <= 0000011101011111;
		weights[3863] <= 1000001100011011;
		weights[3864] <= 0000001111011100;
		weights[3865] <= 0000110110100101;
		weights[3866] <= 0000110111100000;
		weights[3867] <= 0000101001001100;
		weights[3868] <= 0000001101011010;
		weights[3869] <= 1001001111110100;
		weights[3870] <= 1000001010010111;
		weights[3871] <= 0000110111011100;
		weights[3872] <= 0000011111011100;
		weights[3873] <= 0000011111001100;
		weights[3874] <= 0000011110101001;
		weights[3875] <= 1000000110001000;
		weights[3876] <= 1000000010111110;
		weights[3877] <= 1000110010000100;
		weights[3878] <= 1000101101101011;
		weights[3879] <= 1000011000101110;
		weights[3880] <= 1000001001001001;
		weights[3881] <= 0000011111001011;
		weights[3882] <= 0000101010110110;
		weights[3883] <= 0000010011111101;
		weights[3884] <= 1000111100101010;
		weights[3885] <= 0000001011011101;
		weights[3886] <= 1000100111110111;
		weights[3887] <= 1000000010110011;
		weights[3888] <= 1000011001100100;
		weights[3889] <= 1000011010101110;
		weights[3890] <= 0000000001010101;
		weights[3891] <= 0000001000111001;
		weights[3892] <= 1000000011110101;
		weights[3893] <= 0000011000110100;
		weights[3894] <= 0000001100010010;
		weights[3895] <= 0000011010000011;
		weights[3896] <= 0000101111010010;
		weights[3897] <= 1000101001100010;
		weights[3898] <= 1001011000100111;
		weights[3899] <= 1000110111111110;
		weights[3900] <= 1000000101111001;
		weights[3901] <= 0000101010010100;
		weights[3902] <= 0000101110100011;
		weights[3903] <= 0000110110101001;
		weights[3904] <= 1000000101110100;
		weights[3905] <= 1000001100000101;
		weights[3906] <= 1000000110111010;
		weights[3907] <= 0000011100001100;
		weights[3908] <= 0000000001011010;
		weights[3909] <= 1000101110011110;
		weights[3910] <= 0000000011000000;
		weights[3911] <= 1000000111000101;
		weights[3912] <= 0000011100101011;
		weights[3913] <= 1000110011110111;
		weights[3914] <= 0000011111000000;
		weights[3915] <= 1000001110101111;
		weights[3916] <= 0000000111100011;
		weights[3917] <= 0000001000000101;
		weights[3918] <= 1000001110010000;
		weights[3919] <= 0000110100010001;
		weights[3920] <= 0000110001001001;
		weights[3921] <= 0000110100111001;
		weights[3922] <= 1001001001100101;
		weights[3923] <= 1000101000011101;
		weights[3924] <= 1000010101111100;
		weights[3925] <= 0000100011011111;
		weights[3926] <= 1000001000110000;
		weights[3927] <= 1001000100111010;
		weights[3928] <= 1000000010101101;
		weights[3929] <= 1000000111000011;
		weights[3930] <= 0000001000001010;
		weights[3931] <= 1000011000100110;
		weights[3932] <= 0000010000001000;
		weights[3933] <= 1000010001011000;
		weights[3934] <= 1000010110100110;
		weights[3935] <= 0000100110000100;
		weights[3936] <= 0000000000011001;
		weights[3937] <= 1000011010001110;
		weights[3938] <= 1000011110111101;
		weights[3939] <= 0000001110101111;
		weights[3940] <= 1000010101000101;
		weights[3941] <= 1000000111100001;
		weights[3942] <= 0000000000110100;
		weights[3943] <= 1000010110110111;
		weights[3944] <= 1000001100110101;
		weights[3945] <= 1000000011101001;
		weights[3946] <= 1000110001010101;
		weights[3947] <= 0000100011001110;
		weights[3948] <= 1000001101111010;
		weights[3949] <= 1000101101000111;
		weights[3950] <= 0000010011001101;
		weights[3951] <= 0000100000001011;
		weights[3952] <= 0000001111001111;
		weights[3953] <= 1000100100000100;
		weights[3954] <= 1000001110011110;
		weights[3955] <= 1000001011011011;
		weights[3956] <= 0000001110111100;
		weights[3957] <= 1000000010111101;
		weights[3958] <= 1000000011100001;
		weights[3959] <= 0000011101010111;
		weights[3960] <= 1000001100010011;
		weights[3961] <= 0000000110001100;
		weights[3962] <= 1000000010101111;
		weights[3963] <= 0000101001011100;
		weights[3964] <= 0000000111000000;
		weights[3965] <= 0000000110111000;
		weights[3966] <= 0000010110101011;
		weights[3967] <= 0000000011111111;
		weights[3968] <= 1000011101000110;
		weights[3969] <= 1000011001111111;
		weights[3970] <= 1000001010111000;
		weights[3971] <= 0000101011001010;
		weights[3972] <= 1000010100100101;
		weights[3973] <= 1000001010111010;
		weights[3974] <= 1000001001101100;
		weights[3975] <= 0000001101101011;
		weights[3976] <= 1000000111001010;
		weights[3977] <= 1000111000001001;
		weights[3978] <= 1000101101010001;
		weights[3979] <= 0000001100111100;
		weights[3980] <= 1000110101000000;
		weights[3981] <= 0000110001010011;
		weights[3982] <= 0000001010010011;
		weights[3983] <= 0000010011110111;
		weights[3984] <= 1000000001101100;
		weights[3985] <= 1000000111110011;
		weights[3986] <= 1000110011110010;
		weights[3987] <= 0000000011000001;
		weights[3988] <= 1000011000100011;
		weights[3989] <= 0000001101001110;
		weights[3990] <= 0000000100011100;
		weights[3991] <= 0000010101010010;
		weights[3992] <= 1000100000000101;
		weights[3993] <= 1000101000110111;
		weights[3994] <= 1000110001001010;
		weights[3995] <= 0000010110010111;
		weights[3996] <= 0000000110110110;
		weights[3997] <= 0000000100010010;
		weights[3998] <= 1000100010000110;
		weights[3999] <= 0000100000011100;
		weights[4000] <= 1000000100010000;
		weights[4001] <= 0000001111011100;
		weights[4002] <= 0000101000010100;
		weights[4003] <= 0000111000100011;
		weights[4004] <= 1000010100100001;
		weights[4005] <= 0000011100000000;
		weights[4006] <= 0000111100010110;
		weights[4007] <= 0000001001000000;
		weights[4008] <= 0000101110011100;
		weights[4009] <= 0000010001011110;
		weights[4010] <= 1001100011010010;
		weights[4011] <= 0001100100110001;
		weights[4012] <= 1001011001100111;
		weights[4013] <= 1001101010110011;
		weights[4014] <= 0010111010111110;
		weights[4015] <= 0000000001000101;
		weights[4016] <= 0001100100000100;
		weights[4017] <= 0001000010101001;
		weights[4018] <= 1010010000110001;
		weights[4019] <= 0001110000111100;
		weights[4020] <= 1010010110101100;
		weights[4021] <= 1000001011100111;
		weights[4022] <= 0001000001011010;
		weights[4023] <= 0000110000111110;
		weights[4024] <= 1000110110011001;
		weights[4025] <= 0001100111000011;
		weights[4026] <= 0001110101111101;
		weights[4027] <= 1001110111110111;
		weights[4028] <= 1011001110100011;
		weights[4029] <= 1000001101011010;
		weights[4030] <= 1000111010110001;
		weights[4031] <= 1001000110101011;
		weights[4032] <= 1000100100110110;
		weights[4033] <= 0001100101110000;
		weights[4034] <= 1010010000001110;
		weights[4035] <= 0000000011010101;
		weights[4036] <= 1010110110010011;
		weights[4037] <= 0000111000011001;
		weights[4038] <= 1001001100110100;
		weights[4039] <= 0001001000001001;
		weights[4040] <= 1000100011011010;
		weights[4041] <= 0000110110110010;
		weights[4042] <= 0000011101010111;
		weights[4043] <= 0000010000000100;
		weights[4044] <= 1011001000011110;
		weights[4045] <= 0000010100001010;
		weights[4046] <= 0000010100111000;
		weights[4047] <= 1000010110110111;
		weights[4048] <= 1001001101011101;
		weights[4049] <= 1000011001001101;
		weights[4050] <= 0001000011111001;
		weights[4051] <= 0001100000000111;
		weights[4052] <= 0001101110100000;
		weights[4053] <= 1001100011110010;
		weights[4054] <= 1010110100001101;
		weights[4055] <= 0001101010010000;
		weights[4056] <= 0010111011011111;
		weights[4057] <= 1010100001000111;
		weights[4058] <= 0000011101101110;
		weights[4059] <= 1000011101001111;
		weights[4060] <= 0001000101101011;
		weights[4061] <= 0010101111111010;
		weights[4062] <= 0001011011010000;
		weights[4063] <= 1010001100101110;
		weights[4064] <= 1010100011010101;
	end


	always @(negedge(clk)) begin
		if(enable) begin
			case(address)
				12'd0		: data <= weights[0];
				12'd1		: data <= weights[1];
				12'd2		: data <= weights[2];
				12'd3		: data <= weights[3];
				12'd4		: data <= weights[4];
				12'd5		: data <= weights[5];
				12'd6		: data <= weights[6];
				12'd7		: data <= weights[7];
				12'd8		: data <= weights[8];
				12'd9		: data <= weights[9];
				12'd10		: data <= weights[10];
				12'd11		: data <= weights[11];
				12'd12		: data <= weights[12];
				12'd13		: data <= weights[13];
				12'd14		: data <= weights[14];
				12'd15		: data <= weights[15];
				12'd16		: data <= weights[16];
				12'd17		: data <= weights[17];
				12'd18		: data <= weights[18];
				12'd19		: data <= weights[19];
				12'd20		: data <= weights[20];
				12'd21		: data <= weights[21];
				12'd22		: data <= weights[22];
				12'd23		: data <= weights[23];
				12'd24		: data <= weights[24];
				12'd25		: data <= weights[25];
				12'd26		: data <= weights[26];
				12'd27		: data <= weights[27];
				12'd28		: data <= weights[28];
				12'd29		: data <= weights[29];
				12'd30		: data <= weights[30];
				12'd31		: data <= weights[31];
				12'd32		: data <= weights[32];
				12'd33		: data <= weights[33];
				12'd34		: data <= weights[34];
				12'd35		: data <= weights[35];
				12'd36		: data <= weights[36];
				12'd37		: data <= weights[37];
				12'd38		: data <= weights[38];
				12'd39		: data <= weights[39];
				12'd40		: data <= weights[40];
				12'd41		: data <= weights[41];
				12'd42		: data <= weights[42];
				12'd43		: data <= weights[43];
				12'd44		: data <= weights[44];
				12'd45		: data <= weights[45];
				12'd46		: data <= weights[46];
				12'd47		: data <= weights[47];
				12'd48		: data <= weights[48];
				12'd49		: data <= weights[49];
				12'd50		: data <= weights[50];
				12'd51		: data <= weights[51];
				12'd52		: data <= weights[52];
				12'd53		: data <= weights[53];
				12'd54		: data <= weights[54];
				12'd55		: data <= weights[55];
				12'd56		: data <= weights[56];
				12'd57		: data <= weights[57];
				12'd58		: data <= weights[58];
				12'd59		: data <= weights[59];
				12'd60		: data <= weights[60];
				12'd61		: data <= weights[61];
				12'd62		: data <= weights[62];
				12'd63		: data <= weights[63];
				12'd64		: data <= weights[64];
				12'd65		: data <= weights[65];
				12'd66		: data <= weights[66];
				12'd67		: data <= weights[67];
				12'd68		: data <= weights[68];
				12'd69		: data <= weights[69];
				12'd70		: data <= weights[70];
				12'd71		: data <= weights[71];
				12'd72		: data <= weights[72];
				12'd73		: data <= weights[73];
				12'd74		: data <= weights[74];
				12'd75		: data <= weights[75];
				12'd76		: data <= weights[76];
				12'd77		: data <= weights[77];
				12'd78		: data <= weights[78];
				12'd79		: data <= weights[79];
				12'd80		: data <= weights[80];
				12'd81		: data <= weights[81];
				12'd82		: data <= weights[82];
				12'd83		: data <= weights[83];
				12'd84		: data <= weights[84];
				12'd85		: data <= weights[85];
				12'd86		: data <= weights[86];
				12'd87		: data <= weights[87];
				12'd88		: data <= weights[88];
				12'd89		: data <= weights[89];
				12'd90		: data <= weights[90];
				12'd91		: data <= weights[91];
				12'd92		: data <= weights[92];
				12'd93		: data <= weights[93];
				12'd94		: data <= weights[94];
				12'd95		: data <= weights[95];
				12'd96		: data <= weights[96];
				12'd97		: data <= weights[97];
				12'd98		: data <= weights[98];
				12'd99		: data <= weights[99];
				12'd100		: data <= weights[100];
				12'd101		: data <= weights[101];
				12'd102		: data <= weights[102];
				12'd103		: data <= weights[103];
				12'd104		: data <= weights[104];
				12'd105		: data <= weights[105];
				12'd106		: data <= weights[106];
				12'd107		: data <= weights[107];
				12'd108		: data <= weights[108];
				12'd109		: data <= weights[109];
				12'd110		: data <= weights[110];
				12'd111		: data <= weights[111];
				12'd112		: data <= weights[112];
				12'd113		: data <= weights[113];
				12'd114		: data <= weights[114];
				12'd115		: data <= weights[115];
				12'd116		: data <= weights[116];
				12'd117		: data <= weights[117];
				12'd118		: data <= weights[118];
				12'd119		: data <= weights[119];
				12'd120		: data <= weights[120];
				12'd121		: data <= weights[121];
				12'd122		: data <= weights[122];
				12'd123		: data <= weights[123];
				12'd124		: data <= weights[124];
				12'd125		: data <= weights[125];
				12'd126		: data <= weights[126];
				12'd127		: data <= weights[127];
				12'd128		: data <= weights[128];
				12'd129		: data <= weights[129];
				12'd130		: data <= weights[130];
				12'd131		: data <= weights[131];
				12'd132		: data <= weights[132];
				12'd133		: data <= weights[133];
				12'd134		: data <= weights[134];
				12'd135		: data <= weights[135];
				12'd136		: data <= weights[136];
				12'd137		: data <= weights[137];
				12'd138		: data <= weights[138];
				12'd139		: data <= weights[139];
				12'd140		: data <= weights[140];
				12'd141		: data <= weights[141];
				12'd142		: data <= weights[142];
				12'd143		: data <= weights[143];
				12'd144		: data <= weights[144];
				12'd145		: data <= weights[145];
				12'd146		: data <= weights[146];
				12'd147		: data <= weights[147];
				12'd148		: data <= weights[148];
				12'd149		: data <= weights[149];
				12'd150		: data <= weights[150];
				12'd151		: data <= weights[151];
				12'd152		: data <= weights[152];
				12'd153		: data <= weights[153];
				12'd154		: data <= weights[154];
				12'd155		: data <= weights[155];
				12'd156		: data <= weights[156];
				12'd157		: data <= weights[157];
				12'd158		: data <= weights[158];
				12'd159		: data <= weights[159];
				12'd160		: data <= weights[160];
				12'd161		: data <= weights[161];
				12'd162		: data <= weights[162];
				12'd163		: data <= weights[163];
				12'd164		: data <= weights[164];
				12'd165		: data <= weights[165];
				12'd166		: data <= weights[166];
				12'd167		: data <= weights[167];
				12'd168		: data <= weights[168];
				12'd169		: data <= weights[169];
				12'd170		: data <= weights[170];
				12'd171		: data <= weights[171];
				12'd172		: data <= weights[172];
				12'd173		: data <= weights[173];
				12'd174		: data <= weights[174];
				12'd175		: data <= weights[175];
				12'd176		: data <= weights[176];
				12'd177		: data <= weights[177];
				12'd178		: data <= weights[178];
				12'd179		: data <= weights[179];
				12'd180		: data <= weights[180];
				12'd181		: data <= weights[181];
				12'd182		: data <= weights[182];
				12'd183		: data <= weights[183];
				12'd184		: data <= weights[184];
				12'd185		: data <= weights[185];
				12'd186		: data <= weights[186];
				12'd187		: data <= weights[187];
				12'd188		: data <= weights[188];
				12'd189		: data <= weights[189];
				12'd190		: data <= weights[190];
				12'd191		: data <= weights[191];
				12'd192		: data <= weights[192];
				12'd193		: data <= weights[193];
				12'd194		: data <= weights[194];
				12'd195		: data <= weights[195];
				12'd196		: data <= weights[196];
				12'd197		: data <= weights[197];
				12'd198		: data <= weights[198];
				12'd199		: data <= weights[199];
				12'd200		: data <= weights[200];
				12'd201		: data <= weights[201];
				12'd202		: data <= weights[202];
				12'd203		: data <= weights[203];
				12'd204		: data <= weights[204];
				12'd205		: data <= weights[205];
				12'd206		: data <= weights[206];
				12'd207		: data <= weights[207];
				12'd208		: data <= weights[208];
				12'd209		: data <= weights[209];
				12'd210		: data <= weights[210];
				12'd211		: data <= weights[211];
				12'd212		: data <= weights[212];
				12'd213		: data <= weights[213];
				12'd214		: data <= weights[214];
				12'd215		: data <= weights[215];
				12'd216		: data <= weights[216];
				12'd217		: data <= weights[217];
				12'd218		: data <= weights[218];
				12'd219		: data <= weights[219];
				12'd220		: data <= weights[220];
				12'd221		: data <= weights[221];
				12'd222		: data <= weights[222];
				12'd223		: data <= weights[223];
				12'd224		: data <= weights[224];
				12'd225		: data <= weights[225];
				12'd226		: data <= weights[226];
				12'd227		: data <= weights[227];
				12'd228		: data <= weights[228];
				12'd229		: data <= weights[229];
				12'd230		: data <= weights[230];
				12'd231		: data <= weights[231];
				12'd232		: data <= weights[232];
				12'd233		: data <= weights[233];
				12'd234		: data <= weights[234];
				12'd235		: data <= weights[235];
				12'd236		: data <= weights[236];
				12'd237		: data <= weights[237];
				12'd238		: data <= weights[238];
				12'd239		: data <= weights[239];
				12'd240		: data <= weights[240];
				12'd241		: data <= weights[241];
				12'd242		: data <= weights[242];
				12'd243		: data <= weights[243];
				12'd244		: data <= weights[244];
				12'd245		: data <= weights[245];
				12'd246		: data <= weights[246];
				12'd247		: data <= weights[247];
				12'd248		: data <= weights[248];
				12'd249		: data <= weights[249];
				12'd250		: data <= weights[250];
				12'd251		: data <= weights[251];
				12'd252		: data <= weights[252];
				12'd253		: data <= weights[253];
				12'd254		: data <= weights[254];
				12'd255		: data <= weights[255];
				12'd256		: data <= weights[256];
				12'd257		: data <= weights[257];
				12'd258		: data <= weights[258];
				12'd259		: data <= weights[259];
				12'd260		: data <= weights[260];
				12'd261		: data <= weights[261];
				12'd262		: data <= weights[262];
				12'd263		: data <= weights[263];
				12'd264		: data <= weights[264];
				12'd265		: data <= weights[265];
				12'd266		: data <= weights[266];
				12'd267		: data <= weights[267];
				12'd268		: data <= weights[268];
				12'd269		: data <= weights[269];
				12'd270		: data <= weights[270];
				12'd271		: data <= weights[271];
				12'd272		: data <= weights[272];
				12'd273		: data <= weights[273];
				12'd274		: data <= weights[274];
				12'd275		: data <= weights[275];
				12'd276		: data <= weights[276];
				12'd277		: data <= weights[277];
				12'd278		: data <= weights[278];
				12'd279		: data <= weights[279];
				12'd280		: data <= weights[280];
				12'd281		: data <= weights[281];
				12'd282		: data <= weights[282];
				12'd283		: data <= weights[283];
				12'd284		: data <= weights[284];
				12'd285		: data <= weights[285];
				12'd286		: data <= weights[286];
				12'd287		: data <= weights[287];
				12'd288		: data <= weights[288];
				12'd289		: data <= weights[289];
				12'd290		: data <= weights[290];
				12'd291		: data <= weights[291];
				12'd292		: data <= weights[292];
				12'd293		: data <= weights[293];
				12'd294		: data <= weights[294];
				12'd295		: data <= weights[295];
				12'd296		: data <= weights[296];
				12'd297		: data <= weights[297];
				12'd298		: data <= weights[298];
				12'd299		: data <= weights[299];
				12'd300		: data <= weights[300];
				12'd301		: data <= weights[301];
				12'd302		: data <= weights[302];
				12'd303		: data <= weights[303];
				12'd304		: data <= weights[304];
				12'd305		: data <= weights[305];
				12'd306		: data <= weights[306];
				12'd307		: data <= weights[307];
				12'd308		: data <= weights[308];
				12'd309		: data <= weights[309];
				12'd310		: data <= weights[310];
				12'd311		: data <= weights[311];
				12'd312		: data <= weights[312];
				12'd313		: data <= weights[313];
				12'd314		: data <= weights[314];
				12'd315		: data <= weights[315];
				12'd316		: data <= weights[316];
				12'd317		: data <= weights[317];
				12'd318		: data <= weights[318];
				12'd319		: data <= weights[319];
				12'd320		: data <= weights[320];
				12'd321		: data <= weights[321];
				12'd322		: data <= weights[322];
				12'd323		: data <= weights[323];
				12'd324		: data <= weights[324];
				12'd325		: data <= weights[325];
				12'd326		: data <= weights[326];
				12'd327		: data <= weights[327];
				12'd328		: data <= weights[328];
				12'd329		: data <= weights[329];
				12'd330		: data <= weights[330];
				12'd331		: data <= weights[331];
				12'd332		: data <= weights[332];
				12'd333		: data <= weights[333];
				12'd334		: data <= weights[334];
				12'd335		: data <= weights[335];
				12'd336		: data <= weights[336];
				12'd337		: data <= weights[337];
				12'd338		: data <= weights[338];
				12'd339		: data <= weights[339];
				12'd340		: data <= weights[340];
				12'd341		: data <= weights[341];
				12'd342		: data <= weights[342];
				12'd343		: data <= weights[343];
				12'd344		: data <= weights[344];
				12'd345		: data <= weights[345];
				12'd346		: data <= weights[346];
				12'd347		: data <= weights[347];
				12'd348		: data <= weights[348];
				12'd349		: data <= weights[349];
				12'd350		: data <= weights[350];
				12'd351		: data <= weights[351];
				12'd352		: data <= weights[352];
				12'd353		: data <= weights[353];
				12'd354		: data <= weights[354];
				12'd355		: data <= weights[355];
				12'd356		: data <= weights[356];
				12'd357		: data <= weights[357];
				12'd358		: data <= weights[358];
				12'd359		: data <= weights[359];
				12'd360		: data <= weights[360];
				12'd361		: data <= weights[361];
				12'd362		: data <= weights[362];
				12'd363		: data <= weights[363];
				12'd364		: data <= weights[364];
				12'd365		: data <= weights[365];
				12'd366		: data <= weights[366];
				12'd367		: data <= weights[367];
				12'd368		: data <= weights[368];
				12'd369		: data <= weights[369];
				12'd370		: data <= weights[370];
				12'd371		: data <= weights[371];
				12'd372		: data <= weights[372];
				12'd373		: data <= weights[373];
				12'd374		: data <= weights[374];
				12'd375		: data <= weights[375];
				12'd376		: data <= weights[376];
				12'd377		: data <= weights[377];
				12'd378		: data <= weights[378];
				12'd379		: data <= weights[379];
				12'd380		: data <= weights[380];
				12'd381		: data <= weights[381];
				12'd382		: data <= weights[382];
				12'd383		: data <= weights[383];
				12'd384		: data <= weights[384];
				12'd385		: data <= weights[385];
				12'd386		: data <= weights[386];
				12'd387		: data <= weights[387];
				12'd388		: data <= weights[388];
				12'd389		: data <= weights[389];
				12'd390		: data <= weights[390];
				12'd391		: data <= weights[391];
				12'd392		: data <= weights[392];
				12'd393		: data <= weights[393];
				12'd394		: data <= weights[394];
				12'd395		: data <= weights[395];
				12'd396		: data <= weights[396];
				12'd397		: data <= weights[397];
				12'd398		: data <= weights[398];
				12'd399		: data <= weights[399];
				12'd400		: data <= weights[400];
				12'd401		: data <= weights[401];
				12'd402		: data <= weights[402];
				12'd403		: data <= weights[403];
				12'd404		: data <= weights[404];
				12'd405		: data <= weights[405];
				12'd406		: data <= weights[406];
				12'd407		: data <= weights[407];
				12'd408		: data <= weights[408];
				12'd409		: data <= weights[409];
				12'd410		: data <= weights[410];
				12'd411		: data <= weights[411];
				12'd412		: data <= weights[412];
				12'd413		: data <= weights[413];
				12'd414		: data <= weights[414];
				12'd415		: data <= weights[415];
				12'd416		: data <= weights[416];
				12'd417		: data <= weights[417];
				12'd418		: data <= weights[418];
				12'd419		: data <= weights[419];
				12'd420		: data <= weights[420];
				12'd421		: data <= weights[421];
				12'd422		: data <= weights[422];
				12'd423		: data <= weights[423];
				12'd424		: data <= weights[424];
				12'd425		: data <= weights[425];
				12'd426		: data <= weights[426];
				12'd427		: data <= weights[427];
				12'd428		: data <= weights[428];
				12'd429		: data <= weights[429];
				12'd430		: data <= weights[430];
				12'd431		: data <= weights[431];
				12'd432		: data <= weights[432];
				12'd433		: data <= weights[433];
				12'd434		: data <= weights[434];
				12'd435		: data <= weights[435];
				12'd436		: data <= weights[436];
				12'd437		: data <= weights[437];
				12'd438		: data <= weights[438];
				12'd439		: data <= weights[439];
				12'd440		: data <= weights[440];
				12'd441		: data <= weights[441];
				12'd442		: data <= weights[442];
				12'd443		: data <= weights[443];
				12'd444		: data <= weights[444];
				12'd445		: data <= weights[445];
				12'd446		: data <= weights[446];
				12'd447		: data <= weights[447];
				12'd448		: data <= weights[448];
				12'd449		: data <= weights[449];
				12'd450		: data <= weights[450];
				12'd451		: data <= weights[451];
				12'd452		: data <= weights[452];
				12'd453		: data <= weights[453];
				12'd454		: data <= weights[454];
				12'd455		: data <= weights[455];
				12'd456		: data <= weights[456];
				12'd457		: data <= weights[457];
				12'd458		: data <= weights[458];
				12'd459		: data <= weights[459];
				12'd460		: data <= weights[460];
				12'd461		: data <= weights[461];
				12'd462		: data <= weights[462];
				12'd463		: data <= weights[463];
				12'd464		: data <= weights[464];
				12'd465		: data <= weights[465];
				12'd466		: data <= weights[466];
				12'd467		: data <= weights[467];
				12'd468		: data <= weights[468];
				12'd469		: data <= weights[469];
				12'd470		: data <= weights[470];
				12'd471		: data <= weights[471];
				12'd472		: data <= weights[472];
				12'd473		: data <= weights[473];
				12'd474		: data <= weights[474];
				12'd475		: data <= weights[475];
				12'd476		: data <= weights[476];
				12'd477		: data <= weights[477];
				12'd478		: data <= weights[478];
				12'd479		: data <= weights[479];
				12'd480		: data <= weights[480];
				12'd481		: data <= weights[481];
				12'd482		: data <= weights[482];
				12'd483		: data <= weights[483];
				12'd484		: data <= weights[484];
				12'd485		: data <= weights[485];
				12'd486		: data <= weights[486];
				12'd487		: data <= weights[487];
				12'd488		: data <= weights[488];
				12'd489		: data <= weights[489];
				12'd490		: data <= weights[490];
				12'd491		: data <= weights[491];
				12'd492		: data <= weights[492];
				12'd493		: data <= weights[493];
				12'd494		: data <= weights[494];
				12'd495		: data <= weights[495];
				12'd496		: data <= weights[496];
				12'd497		: data <= weights[497];
				12'd498		: data <= weights[498];
				12'd499		: data <= weights[499];
				12'd500		: data <= weights[500];
				12'd501		: data <= weights[501];
				12'd502		: data <= weights[502];
				12'd503		: data <= weights[503];
				12'd504		: data <= weights[504];
				12'd505		: data <= weights[505];
				12'd506		: data <= weights[506];
				12'd507		: data <= weights[507];
				12'd508		: data <= weights[508];
				12'd509		: data <= weights[509];
				12'd510		: data <= weights[510];
				12'd511		: data <= weights[511];
				12'd512		: data <= weights[512];
				12'd513		: data <= weights[513];
				12'd514		: data <= weights[514];
				12'd515		: data <= weights[515];
				12'd516		: data <= weights[516];
				12'd517		: data <= weights[517];
				12'd518		: data <= weights[518];
				12'd519		: data <= weights[519];
				12'd520		: data <= weights[520];
				12'd521		: data <= weights[521];
				12'd522		: data <= weights[522];
				12'd523		: data <= weights[523];
				12'd524		: data <= weights[524];
				12'd525		: data <= weights[525];
				12'd526		: data <= weights[526];
				12'd527		: data <= weights[527];
				12'd528		: data <= weights[528];
				12'd529		: data <= weights[529];
				12'd530		: data <= weights[530];
				12'd531		: data <= weights[531];
				12'd532		: data <= weights[532];
				12'd533		: data <= weights[533];
				12'd534		: data <= weights[534];
				12'd535		: data <= weights[535];
				12'd536		: data <= weights[536];
				12'd537		: data <= weights[537];
				12'd538		: data <= weights[538];
				12'd539		: data <= weights[539];
				12'd540		: data <= weights[540];
				12'd541		: data <= weights[541];
				12'd542		: data <= weights[542];
				12'd543		: data <= weights[543];
				12'd544		: data <= weights[544];
				12'd545		: data <= weights[545];
				12'd546		: data <= weights[546];
				12'd547		: data <= weights[547];
				12'd548		: data <= weights[548];
				12'd549		: data <= weights[549];
				12'd550		: data <= weights[550];
				12'd551		: data <= weights[551];
				12'd552		: data <= weights[552];
				12'd553		: data <= weights[553];
				12'd554		: data <= weights[554];
				12'd555		: data <= weights[555];
				12'd556		: data <= weights[556];
				12'd557		: data <= weights[557];
				12'd558		: data <= weights[558];
				12'd559		: data <= weights[559];
				12'd560		: data <= weights[560];
				12'd561		: data <= weights[561];
				12'd562		: data <= weights[562];
				12'd563		: data <= weights[563];
				12'd564		: data <= weights[564];
				12'd565		: data <= weights[565];
				12'd566		: data <= weights[566];
				12'd567		: data <= weights[567];
				12'd568		: data <= weights[568];
				12'd569		: data <= weights[569];
				12'd570		: data <= weights[570];
				12'd571		: data <= weights[571];
				12'd572		: data <= weights[572];
				12'd573		: data <= weights[573];
				12'd574		: data <= weights[574];
				12'd575		: data <= weights[575];
				12'd576		: data <= weights[576];
				12'd577		: data <= weights[577];
				12'd578		: data <= weights[578];
				12'd579		: data <= weights[579];
				12'd580		: data <= weights[580];
				12'd581		: data <= weights[581];
				12'd582		: data <= weights[582];
				12'd583		: data <= weights[583];
				12'd584		: data <= weights[584];
				12'd585		: data <= weights[585];
				12'd586		: data <= weights[586];
				12'd587		: data <= weights[587];
				12'd588		: data <= weights[588];
				12'd589		: data <= weights[589];
				12'd590		: data <= weights[590];
				12'd591		: data <= weights[591];
				12'd592		: data <= weights[592];
				12'd593		: data <= weights[593];
				12'd594		: data <= weights[594];
				12'd595		: data <= weights[595];
				12'd596		: data <= weights[596];
				12'd597		: data <= weights[597];
				12'd598		: data <= weights[598];
				12'd599		: data <= weights[599];
				12'd600		: data <= weights[600];
				12'd601		: data <= weights[601];
				12'd602		: data <= weights[602];
				12'd603		: data <= weights[603];
				12'd604		: data <= weights[604];
				12'd605		: data <= weights[605];
				12'd606		: data <= weights[606];
				12'd607		: data <= weights[607];
				12'd608		: data <= weights[608];
				12'd609		: data <= weights[609];
				12'd610		: data <= weights[610];
				12'd611		: data <= weights[611];
				12'd612		: data <= weights[612];
				12'd613		: data <= weights[613];
				12'd614		: data <= weights[614];
				12'd615		: data <= weights[615];
				12'd616		: data <= weights[616];
				12'd617		: data <= weights[617];
				12'd618		: data <= weights[618];
				12'd619		: data <= weights[619];
				12'd620		: data <= weights[620];
				12'd621		: data <= weights[621];
				12'd622		: data <= weights[622];
				12'd623		: data <= weights[623];
				12'd624		: data <= weights[624];
				12'd625		: data <= weights[625];
				12'd626		: data <= weights[626];
				12'd627		: data <= weights[627];
				12'd628		: data <= weights[628];
				12'd629		: data <= weights[629];
				12'd630		: data <= weights[630];
				12'd631		: data <= weights[631];
				12'd632		: data <= weights[632];
				12'd633		: data <= weights[633];
				12'd634		: data <= weights[634];
				12'd635		: data <= weights[635];
				12'd636		: data <= weights[636];
				12'd637		: data <= weights[637];
				12'd638		: data <= weights[638];
				12'd639		: data <= weights[639];
				12'd640		: data <= weights[640];
				12'd641		: data <= weights[641];
				12'd642		: data <= weights[642];
				12'd643		: data <= weights[643];
				12'd644		: data <= weights[644];
				12'd645		: data <= weights[645];
				12'd646		: data <= weights[646];
				12'd647		: data <= weights[647];
				12'd648		: data <= weights[648];
				12'd649		: data <= weights[649];
				12'd650		: data <= weights[650];
				12'd651		: data <= weights[651];
				12'd652		: data <= weights[652];
				12'd653		: data <= weights[653];
				12'd654		: data <= weights[654];
				12'd655		: data <= weights[655];
				12'd656		: data <= weights[656];
				12'd657		: data <= weights[657];
				12'd658		: data <= weights[658];
				12'd659		: data <= weights[659];
				12'd660		: data <= weights[660];
				12'd661		: data <= weights[661];
				12'd662		: data <= weights[662];
				12'd663		: data <= weights[663];
				12'd664		: data <= weights[664];
				12'd665		: data <= weights[665];
				12'd666		: data <= weights[666];
				12'd667		: data <= weights[667];
				12'd668		: data <= weights[668];
				12'd669		: data <= weights[669];
				12'd670		: data <= weights[670];
				12'd671		: data <= weights[671];
				12'd672		: data <= weights[672];
				12'd673		: data <= weights[673];
				12'd674		: data <= weights[674];
				12'd675		: data <= weights[675];
				12'd676		: data <= weights[676];
				12'd677		: data <= weights[677];
				12'd678		: data <= weights[678];
				12'd679		: data <= weights[679];
				12'd680		: data <= weights[680];
				12'd681		: data <= weights[681];
				12'd682		: data <= weights[682];
				12'd683		: data <= weights[683];
				12'd684		: data <= weights[684];
				12'd685		: data <= weights[685];
				12'd686		: data <= weights[686];
				12'd687		: data <= weights[687];
				12'd688		: data <= weights[688];
				12'd689		: data <= weights[689];
				12'd690		: data <= weights[690];
				12'd691		: data <= weights[691];
				12'd692		: data <= weights[692];
				12'd693		: data <= weights[693];
				12'd694		: data <= weights[694];
				12'd695		: data <= weights[695];
				12'd696		: data <= weights[696];
				12'd697		: data <= weights[697];
				12'd698		: data <= weights[698];
				12'd699		: data <= weights[699];
				12'd700		: data <= weights[700];
				12'd701		: data <= weights[701];
				12'd702		: data <= weights[702];
				12'd703		: data <= weights[703];
				12'd704		: data <= weights[704];
				12'd705		: data <= weights[705];
				12'd706		: data <= weights[706];
				12'd707		: data <= weights[707];
				12'd708		: data <= weights[708];
				12'd709		: data <= weights[709];
				12'd710		: data <= weights[710];
				12'd711		: data <= weights[711];
				12'd712		: data <= weights[712];
				12'd713		: data <= weights[713];
				12'd714		: data <= weights[714];
				12'd715		: data <= weights[715];
				12'd716		: data <= weights[716];
				12'd717		: data <= weights[717];
				12'd718		: data <= weights[718];
				12'd719		: data <= weights[719];
				12'd720		: data <= weights[720];
				12'd721		: data <= weights[721];
				12'd722		: data <= weights[722];
				12'd723		: data <= weights[723];
				12'd724		: data <= weights[724];
				12'd725		: data <= weights[725];
				12'd726		: data <= weights[726];
				12'd727		: data <= weights[727];
				12'd728		: data <= weights[728];
				12'd729		: data <= weights[729];
				12'd730		: data <= weights[730];
				12'd731		: data <= weights[731];
				12'd732		: data <= weights[732];
				12'd733		: data <= weights[733];
				12'd734		: data <= weights[734];
				12'd735		: data <= weights[735];
				12'd736		: data <= weights[736];
				12'd737		: data <= weights[737];
				12'd738		: data <= weights[738];
				12'd739		: data <= weights[739];
				12'd740		: data <= weights[740];
				12'd741		: data <= weights[741];
				12'd742		: data <= weights[742];
				12'd743		: data <= weights[743];
				12'd744		: data <= weights[744];
				12'd745		: data <= weights[745];
				12'd746		: data <= weights[746];
				12'd747		: data <= weights[747];
				12'd748		: data <= weights[748];
				12'd749		: data <= weights[749];
				12'd750		: data <= weights[750];
				12'd751		: data <= weights[751];
				12'd752		: data <= weights[752];
				12'd753		: data <= weights[753];
				12'd754		: data <= weights[754];
				12'd755		: data <= weights[755];
				12'd756		: data <= weights[756];
				12'd757		: data <= weights[757];
				12'd758		: data <= weights[758];
				12'd759		: data <= weights[759];
				12'd760		: data <= weights[760];
				12'd761		: data <= weights[761];
				12'd762		: data <= weights[762];
				12'd763		: data <= weights[763];
				12'd764		: data <= weights[764];
				12'd765		: data <= weights[765];
				12'd766		: data <= weights[766];
				12'd767		: data <= weights[767];
				12'd768		: data <= weights[768];
				12'd769		: data <= weights[769];
				12'd770		: data <= weights[770];
				12'd771		: data <= weights[771];
				12'd772		: data <= weights[772];
				12'd773		: data <= weights[773];
				12'd774		: data <= weights[774];
				12'd775		: data <= weights[775];
				12'd776		: data <= weights[776];
				12'd777		: data <= weights[777];
				12'd778		: data <= weights[778];
				12'd779		: data <= weights[779];
				12'd780		: data <= weights[780];
				12'd781		: data <= weights[781];
				12'd782		: data <= weights[782];
				12'd783		: data <= weights[783];
				12'd784		: data <= weights[784];
				12'd785		: data <= weights[785];
				12'd786		: data <= weights[786];
				12'd787		: data <= weights[787];
				12'd788		: data <= weights[788];
				12'd789		: data <= weights[789];
				12'd790		: data <= weights[790];
				12'd791		: data <= weights[791];
				12'd792		: data <= weights[792];
				12'd793		: data <= weights[793];
				12'd794		: data <= weights[794];
				12'd795		: data <= weights[795];
				12'd796		: data <= weights[796];
				12'd797		: data <= weights[797];
				12'd798		: data <= weights[798];
				12'd799		: data <= weights[799];
				12'd800		: data <= weights[800];
				12'd801		: data <= weights[801];
				12'd802		: data <= weights[802];
				12'd803		: data <= weights[803];
				12'd804		: data <= weights[804];
				12'd805		: data <= weights[805];
				12'd806		: data <= weights[806];
				12'd807		: data <= weights[807];
				12'd808		: data <= weights[808];
				12'd809		: data <= weights[809];
				12'd810		: data <= weights[810];
				12'd811		: data <= weights[811];
				12'd812		: data <= weights[812];
				12'd813		: data <= weights[813];
				12'd814		: data <= weights[814];
				12'd815		: data <= weights[815];
				12'd816		: data <= weights[816];
				12'd817		: data <= weights[817];
				12'd818		: data <= weights[818];
				12'd819		: data <= weights[819];
				12'd820		: data <= weights[820];
				12'd821		: data <= weights[821];
				12'd822		: data <= weights[822];
				12'd823		: data <= weights[823];
				12'd824		: data <= weights[824];
				12'd825		: data <= weights[825];
				12'd826		: data <= weights[826];
				12'd827		: data <= weights[827];
				12'd828		: data <= weights[828];
				12'd829		: data <= weights[829];
				12'd830		: data <= weights[830];
				12'd831		: data <= weights[831];
				12'd832		: data <= weights[832];
				12'd833		: data <= weights[833];
				12'd834		: data <= weights[834];
				12'd835		: data <= weights[835];
				12'd836		: data <= weights[836];
				12'd837		: data <= weights[837];
				12'd838		: data <= weights[838];
				12'd839		: data <= weights[839];
				12'd840		: data <= weights[840];
				12'd841		: data <= weights[841];
				12'd842		: data <= weights[842];
				12'd843		: data <= weights[843];
				12'd844		: data <= weights[844];
				12'd845		: data <= weights[845];
				12'd846		: data <= weights[846];
				12'd847		: data <= weights[847];
				12'd848		: data <= weights[848];
				12'd849		: data <= weights[849];
				12'd850		: data <= weights[850];
				12'd851		: data <= weights[851];
				12'd852		: data <= weights[852];
				12'd853		: data <= weights[853];
				12'd854		: data <= weights[854];
				12'd855		: data <= weights[855];
				12'd856		: data <= weights[856];
				12'd857		: data <= weights[857];
				12'd858		: data <= weights[858];
				12'd859		: data <= weights[859];
				12'd860		: data <= weights[860];
				12'd861		: data <= weights[861];
				12'd862		: data <= weights[862];
				12'd863		: data <= weights[863];
				12'd864		: data <= weights[864];
				12'd865		: data <= weights[865];
				12'd866		: data <= weights[866];
				12'd867		: data <= weights[867];
				12'd868		: data <= weights[868];
				12'd869		: data <= weights[869];
				12'd870		: data <= weights[870];
				12'd871		: data <= weights[871];
				12'd872		: data <= weights[872];
				12'd873		: data <= weights[873];
				12'd874		: data <= weights[874];
				12'd875		: data <= weights[875];
				12'd876		: data <= weights[876];
				12'd877		: data <= weights[877];
				12'd878		: data <= weights[878];
				12'd879		: data <= weights[879];
				12'd880		: data <= weights[880];
				12'd881		: data <= weights[881];
				12'd882		: data <= weights[882];
				12'd883		: data <= weights[883];
				12'd884		: data <= weights[884];
				12'd885		: data <= weights[885];
				12'd886		: data <= weights[886];
				12'd887		: data <= weights[887];
				12'd888		: data <= weights[888];
				12'd889		: data <= weights[889];
				12'd890		: data <= weights[890];
				12'd891		: data <= weights[891];
				12'd892		: data <= weights[892];
				12'd893		: data <= weights[893];
				12'd894		: data <= weights[894];
				12'd895		: data <= weights[895];
				12'd896		: data <= weights[896];
				12'd897		: data <= weights[897];
				12'd898		: data <= weights[898];
				12'd899		: data <= weights[899];
				12'd900		: data <= weights[900];
				12'd901		: data <= weights[901];
				12'd902		: data <= weights[902];
				12'd903		: data <= weights[903];
				12'd904		: data <= weights[904];
				12'd905		: data <= weights[905];
				12'd906		: data <= weights[906];
				12'd907		: data <= weights[907];
				12'd908		: data <= weights[908];
				12'd909		: data <= weights[909];
				12'd910		: data <= weights[910];
				12'd911		: data <= weights[911];
				12'd912		: data <= weights[912];
				12'd913		: data <= weights[913];
				12'd914		: data <= weights[914];
				12'd915		: data <= weights[915];
				12'd916		: data <= weights[916];
				12'd917		: data <= weights[917];
				12'd918		: data <= weights[918];
				12'd919		: data <= weights[919];
				12'd920		: data <= weights[920];
				12'd921		: data <= weights[921];
				12'd922		: data <= weights[922];
				12'd923		: data <= weights[923];
				12'd924		: data <= weights[924];
				12'd925		: data <= weights[925];
				12'd926		: data <= weights[926];
				12'd927		: data <= weights[927];
				12'd928		: data <= weights[928];
				12'd929		: data <= weights[929];
				12'd930		: data <= weights[930];
				12'd931		: data <= weights[931];
				12'd932		: data <= weights[932];
				12'd933		: data <= weights[933];
				12'd934		: data <= weights[934];
				12'd935		: data <= weights[935];
				12'd936		: data <= weights[936];
				12'd937		: data <= weights[937];
				12'd938		: data <= weights[938];
				12'd939		: data <= weights[939];
				12'd940		: data <= weights[940];
				12'd941		: data <= weights[941];
				12'd942		: data <= weights[942];
				12'd943		: data <= weights[943];
				12'd944		: data <= weights[944];
				12'd945		: data <= weights[945];
				12'd946		: data <= weights[946];
				12'd947		: data <= weights[947];
				12'd948		: data <= weights[948];
				12'd949		: data <= weights[949];
				12'd950		: data <= weights[950];
				12'd951		: data <= weights[951];
				12'd952		: data <= weights[952];
				12'd953		: data <= weights[953];
				12'd954		: data <= weights[954];
				12'd955		: data <= weights[955];
				12'd956		: data <= weights[956];
				12'd957		: data <= weights[957];
				12'd958		: data <= weights[958];
				12'd959		: data <= weights[959];
				12'd960		: data <= weights[960];
				12'd961		: data <= weights[961];
				12'd962		: data <= weights[962];
				12'd963		: data <= weights[963];
				12'd964		: data <= weights[964];
				12'd965		: data <= weights[965];
				12'd966		: data <= weights[966];
				12'd967		: data <= weights[967];
				12'd968		: data <= weights[968];
				12'd969		: data <= weights[969];
				12'd970		: data <= weights[970];
				12'd971		: data <= weights[971];
				12'd972		: data <= weights[972];
				12'd973		: data <= weights[973];
				12'd974		: data <= weights[974];
				12'd975		: data <= weights[975];
				12'd976		: data <= weights[976];
				12'd977		: data <= weights[977];
				12'd978		: data <= weights[978];
				12'd979		: data <= weights[979];
				12'd980		: data <= weights[980];
				12'd981		: data <= weights[981];
				12'd982		: data <= weights[982];
				12'd983		: data <= weights[983];
				12'd984		: data <= weights[984];
				12'd985		: data <= weights[985];
				12'd986		: data <= weights[986];
				12'd987		: data <= weights[987];
				12'd988		: data <= weights[988];
				12'd989		: data <= weights[989];
				12'd990		: data <= weights[990];
				12'd991		: data <= weights[991];
				12'd992		: data <= weights[992];
				12'd993		: data <= weights[993];
				12'd994		: data <= weights[994];
				12'd995		: data <= weights[995];
				12'd996		: data <= weights[996];
				12'd997		: data <= weights[997];
				12'd998		: data <= weights[998];
				12'd999		: data <= weights[999];
				12'd1000	: data <= weights[1000];
				12'd1001	: data <= weights[1001];
				12'd1002	: data <= weights[1002];
				12'd1003	: data <= weights[1003];
				12'd1004	: data <= weights[1004];
				12'd1005	: data <= weights[1005];
				12'd1006	: data <= weights[1006];
				12'd1007	: data <= weights[1007];
				12'd1008	: data <= weights[1008];
				12'd1009	: data <= weights[1009];
				12'd1010	: data <= weights[1010];
				12'd1011	: data <= weights[1011];
				12'd1012	: data <= weights[1012];
				12'd1013	: data <= weights[1013];
				12'd1014	: data <= weights[1014];
				12'd1015	: data <= weights[1015];
				12'd1016	: data <= weights[1016];
				12'd1017	: data <= weights[1017];
				12'd1018	: data <= weights[1018];
				12'd1019	: data <= weights[1019];
				12'd1020	: data <= weights[1020];
				12'd1021	: data <= weights[1021];
				12'd1022	: data <= weights[1022];
				12'd1023	: data <= weights[1023];
				12'd1024	: data <= weights[1024];
				12'd1025	: data <= weights[1025];
				12'd1026	: data <= weights[1026];
				12'd1027	: data <= weights[1027];
				12'd1028	: data <= weights[1028];
				12'd1029	: data <= weights[1029];
				12'd1030	: data <= weights[1030];
				12'd1031	: data <= weights[1031];
				12'd1032	: data <= weights[1032];
				12'd1033	: data <= weights[1033];
				12'd1034	: data <= weights[1034];
				12'd1035	: data <= weights[1035];
				12'd1036	: data <= weights[1036];
				12'd1037	: data <= weights[1037];
				12'd1038	: data <= weights[1038];
				12'd1039	: data <= weights[1039];
				12'd1040	: data <= weights[1040];
				12'd1041	: data <= weights[1041];
				12'd1042	: data <= weights[1042];
				12'd1043	: data <= weights[1043];
				12'd1044	: data <= weights[1044];
				12'd1045	: data <= weights[1045];
				12'd1046	: data <= weights[1046];
				12'd1047	: data <= weights[1047];
				12'd1048	: data <= weights[1048];
				12'd1049	: data <= weights[1049];
				12'd1050	: data <= weights[1050];
				12'd1051	: data <= weights[1051];
				12'd1052	: data <= weights[1052];
				12'd1053	: data <= weights[1053];
				12'd1054	: data <= weights[1054];
				12'd1055	: data <= weights[1055];
				12'd1056	: data <= weights[1056];
				12'd1057	: data <= weights[1057];
				12'd1058	: data <= weights[1058];
				12'd1059	: data <= weights[1059];
				12'd1060	: data <= weights[1060];
				12'd1061	: data <= weights[1061];
				12'd1062	: data <= weights[1062];
				12'd1063	: data <= weights[1063];
				12'd1064	: data <= weights[1064];
				12'd1065	: data <= weights[1065];
				12'd1066	: data <= weights[1066];
				12'd1067	: data <= weights[1067];
				12'd1068	: data <= weights[1068];
				12'd1069	: data <= weights[1069];
				12'd1070	: data <= weights[1070];
				12'd1071	: data <= weights[1071];
				12'd1072	: data <= weights[1072];
				12'd1073	: data <= weights[1073];
				12'd1074	: data <= weights[1074];
				12'd1075	: data <= weights[1075];
				12'd1076	: data <= weights[1076];
				12'd1077	: data <= weights[1077];
				12'd1078	: data <= weights[1078];
				12'd1079	: data <= weights[1079];
				12'd1080	: data <= weights[1080];
				12'd1081	: data <= weights[1081];
				12'd1082	: data <= weights[1082];
				12'd1083	: data <= weights[1083];
				12'd1084	: data <= weights[1084];
				12'd1085	: data <= weights[1085];
				12'd1086	: data <= weights[1086];
				12'd1087	: data <= weights[1087];
				12'd1088	: data <= weights[1088];
				12'd1089	: data <= weights[1089];
				12'd1090	: data <= weights[1090];
				12'd1091	: data <= weights[1091];
				12'd1092	: data <= weights[1092];
				12'd1093	: data <= weights[1093];
				12'd1094	: data <= weights[1094];
				12'd1095	: data <= weights[1095];
				12'd1096	: data <= weights[1096];
				12'd1097	: data <= weights[1097];
				12'd1098	: data <= weights[1098];
				12'd1099	: data <= weights[1099];
				12'd1100	: data <= weights[1100];
				12'd1101	: data <= weights[1101];
				12'd1102	: data <= weights[1102];
				12'd1103	: data <= weights[1103];
				12'd1104	: data <= weights[1104];
				12'd1105	: data <= weights[1105];
				12'd1106	: data <= weights[1106];
				12'd1107	: data <= weights[1107];
				12'd1108	: data <= weights[1108];
				12'd1109	: data <= weights[1109];
				12'd1110	: data <= weights[1110];
				12'd1111	: data <= weights[1111];
				12'd1112	: data <= weights[1112];
				12'd1113	: data <= weights[1113];
				12'd1114	: data <= weights[1114];
				12'd1115	: data <= weights[1115];
				12'd1116	: data <= weights[1116];
				12'd1117	: data <= weights[1117];
				12'd1118	: data <= weights[1118];
				12'd1119	: data <= weights[1119];
				12'd1120	: data <= weights[1120];
				12'd1121	: data <= weights[1121];
				12'd1122	: data <= weights[1122];
				12'd1123	: data <= weights[1123];
				12'd1124	: data <= weights[1124];
				12'd1125	: data <= weights[1125];
				12'd1126	: data <= weights[1126];
				12'd1127	: data <= weights[1127];
				12'd1128	: data <= weights[1128];
				12'd1129	: data <= weights[1129];
				12'd1130	: data <= weights[1130];
				12'd1131	: data <= weights[1131];
				12'd1132	: data <= weights[1132];
				12'd1133	: data <= weights[1133];
				12'd1134	: data <= weights[1134];
				12'd1135	: data <= weights[1135];
				12'd1136	: data <= weights[1136];
				12'd1137	: data <= weights[1137];
				12'd1138	: data <= weights[1138];
				12'd1139	: data <= weights[1139];
				12'd1140	: data <= weights[1140];
				12'd1141	: data <= weights[1141];
				12'd1142	: data <= weights[1142];
				12'd1143	: data <= weights[1143];
				12'd1144	: data <= weights[1144];
				12'd1145	: data <= weights[1145];
				12'd1146	: data <= weights[1146];
				12'd1147	: data <= weights[1147];
				12'd1148	: data <= weights[1148];
				12'd1149	: data <= weights[1149];
				12'd1150	: data <= weights[1150];
				12'd1151	: data <= weights[1151];
				12'd1152	: data <= weights[1152];
				12'd1153	: data <= weights[1153];
				12'd1154	: data <= weights[1154];
				12'd1155	: data <= weights[1155];
				12'd1156	: data <= weights[1156];
				12'd1157	: data <= weights[1157];
				12'd1158	: data <= weights[1158];
				12'd1159	: data <= weights[1159];
				12'd1160	: data <= weights[1160];
				12'd1161	: data <= weights[1161];
				12'd1162	: data <= weights[1162];
				12'd1163	: data <= weights[1163];
				12'd1164	: data <= weights[1164];
				12'd1165	: data <= weights[1165];
				12'd1166	: data <= weights[1166];
				12'd1167	: data <= weights[1167];
				12'd1168	: data <= weights[1168];
				12'd1169	: data <= weights[1169];
				12'd1170	: data <= weights[1170];
				12'd1171	: data <= weights[1171];
				12'd1172	: data <= weights[1172];
				12'd1173	: data <= weights[1173];
				12'd1174	: data <= weights[1174];
				12'd1175	: data <= weights[1175];
				12'd1176	: data <= weights[1176];
				12'd1177	: data <= weights[1177];
				12'd1178	: data <= weights[1178];
				12'd1179	: data <= weights[1179];
				12'd1180	: data <= weights[1180];
				12'd1181	: data <= weights[1181];
				12'd1182	: data <= weights[1182];
				12'd1183	: data <= weights[1183];
				12'd1184	: data <= weights[1184];
				12'd1185	: data <= weights[1185];
				12'd1186	: data <= weights[1186];
				12'd1187	: data <= weights[1187];
				12'd1188	: data <= weights[1188];
				12'd1189	: data <= weights[1189];
				12'd1190	: data <= weights[1190];
				12'd1191	: data <= weights[1191];
				12'd1192	: data <= weights[1192];
				12'd1193	: data <= weights[1193];
				12'd1194	: data <= weights[1194];
				12'd1195	: data <= weights[1195];
				12'd1196	: data <= weights[1196];
				12'd1197	: data <= weights[1197];
				12'd1198	: data <= weights[1198];
				12'd1199	: data <= weights[1199];
				12'd1200	: data <= weights[1200];
				12'd1201	: data <= weights[1201];
				12'd1202	: data <= weights[1202];
				12'd1203	: data <= weights[1203];
				12'd1204	: data <= weights[1204];
				12'd1205	: data <= weights[1205];
				12'd1206	: data <= weights[1206];
				12'd1207	: data <= weights[1207];
				12'd1208	: data <= weights[1208];
				12'd1209	: data <= weights[1209];
				12'd1210	: data <= weights[1210];
				12'd1211	: data <= weights[1211];
				12'd1212	: data <= weights[1212];
				12'd1213	: data <= weights[1213];
				12'd1214	: data <= weights[1214];
				12'd1215	: data <= weights[1215];
				12'd1216	: data <= weights[1216];
				12'd1217	: data <= weights[1217];
				12'd1218	: data <= weights[1218];
				12'd1219	: data <= weights[1219];
				12'd1220	: data <= weights[1220];
				12'd1221	: data <= weights[1221];
				12'd1222	: data <= weights[1222];
				12'd1223	: data <= weights[1223];
				12'd1224	: data <= weights[1224];
				12'd1225	: data <= weights[1225];
				12'd1226	: data <= weights[1226];
				12'd1227	: data <= weights[1227];
				12'd1228	: data <= weights[1228];
				12'd1229	: data <= weights[1229];
				12'd1230	: data <= weights[1230];
				12'd1231	: data <= weights[1231];
				12'd1232	: data <= weights[1232];
				12'd1233	: data <= weights[1233];
				12'd1234	: data <= weights[1234];
				12'd1235	: data <= weights[1235];
				12'd1236	: data <= weights[1236];
				12'd1237	: data <= weights[1237];
				12'd1238	: data <= weights[1238];
				12'd1239	: data <= weights[1239];
				12'd1240	: data <= weights[1240];
				12'd1241	: data <= weights[1241];
				12'd1242	: data <= weights[1242];
				12'd1243	: data <= weights[1243];
				12'd1244	: data <= weights[1244];
				12'd1245	: data <= weights[1245];
				12'd1246	: data <= weights[1246];
				12'd1247	: data <= weights[1247];
				12'd1248	: data <= weights[1248];
				12'd1249	: data <= weights[1249];
				12'd1250	: data <= weights[1250];
				12'd1251	: data <= weights[1251];
				12'd1252	: data <= weights[1252];
				12'd1253	: data <= weights[1253];
				12'd1254	: data <= weights[1254];
				12'd1255	: data <= weights[1255];
				12'd1256	: data <= weights[1256];
				12'd1257	: data <= weights[1257];
				12'd1258	: data <= weights[1258];
				12'd1259	: data <= weights[1259];
				12'd1260	: data <= weights[1260];
				12'd1261	: data <= weights[1261];
				12'd1262	: data <= weights[1262];
				12'd1263	: data <= weights[1263];
				12'd1264	: data <= weights[1264];
				12'd1265	: data <= weights[1265];
				12'd1266	: data <= weights[1266];
				12'd1267	: data <= weights[1267];
				12'd1268	: data <= weights[1268];
				12'd1269	: data <= weights[1269];
				12'd1270	: data <= weights[1270];
				12'd1271	: data <= weights[1271];
				12'd1272	: data <= weights[1272];
				12'd1273	: data <= weights[1273];
				12'd1274	: data <= weights[1274];
				12'd1275	: data <= weights[1275];
				12'd1276	: data <= weights[1276];
				12'd1277	: data <= weights[1277];
				12'd1278	: data <= weights[1278];
				12'd1279	: data <= weights[1279];
				12'd1280	: data <= weights[1280];
				12'd1281	: data <= weights[1281];
				12'd1282	: data <= weights[1282];
				12'd1283	: data <= weights[1283];
				12'd1284	: data <= weights[1284];
				12'd1285	: data <= weights[1285];
				12'd1286	: data <= weights[1286];
				12'd1287	: data <= weights[1287];
				12'd1288	: data <= weights[1288];
				12'd1289	: data <= weights[1289];
				12'd1290	: data <= weights[1290];
				12'd1291	: data <= weights[1291];
				12'd1292	: data <= weights[1292];
				12'd1293	: data <= weights[1293];
				12'd1294	: data <= weights[1294];
				12'd1295	: data <= weights[1295];
				12'd1296	: data <= weights[1296];
				12'd1297	: data <= weights[1297];
				12'd1298	: data <= weights[1298];
				12'd1299	: data <= weights[1299];
				12'd1300	: data <= weights[1300];
				12'd1301	: data <= weights[1301];
				12'd1302	: data <= weights[1302];
				12'd1303	: data <= weights[1303];
				12'd1304	: data <= weights[1304];
				12'd1305	: data <= weights[1305];
				12'd1306	: data <= weights[1306];
				12'd1307	: data <= weights[1307];
				12'd1308	: data <= weights[1308];
				12'd1309	: data <= weights[1309];
				12'd1310	: data <= weights[1310];
				12'd1311	: data <= weights[1311];
				12'd1312	: data <= weights[1312];
				12'd1313	: data <= weights[1313];
				12'd1314	: data <= weights[1314];
				12'd1315	: data <= weights[1315];
				12'd1316	: data <= weights[1316];
				12'd1317	: data <= weights[1317];
				12'd1318	: data <= weights[1318];
				12'd1319	: data <= weights[1319];
				12'd1320	: data <= weights[1320];
				12'd1321	: data <= weights[1321];
				12'd1322	: data <= weights[1322];
				12'd1323	: data <= weights[1323];
				12'd1324	: data <= weights[1324];
				12'd1325	: data <= weights[1325];
				12'd1326	: data <= weights[1326];
				12'd1327	: data <= weights[1327];
				12'd1328	: data <= weights[1328];
				12'd1329	: data <= weights[1329];
				12'd1330	: data <= weights[1330];
				12'd1331	: data <= weights[1331];
				12'd1332	: data <= weights[1332];
				12'd1333	: data <= weights[1333];
				12'd1334	: data <= weights[1334];
				12'd1335	: data <= weights[1335];
				12'd1336	: data <= weights[1336];
				12'd1337	: data <= weights[1337];
				12'd1338	: data <= weights[1338];
				12'd1339	: data <= weights[1339];
				12'd1340	: data <= weights[1340];
				12'd1341	: data <= weights[1341];
				12'd1342	: data <= weights[1342];
				12'd1343	: data <= weights[1343];
				12'd1344	: data <= weights[1344];
				12'd1345	: data <= weights[1345];
				12'd1346	: data <= weights[1346];
				12'd1347	: data <= weights[1347];
				12'd1348	: data <= weights[1348];
				12'd1349	: data <= weights[1349];
				12'd1350	: data <= weights[1350];
				12'd1351	: data <= weights[1351];
				12'd1352	: data <= weights[1352];
				12'd1353	: data <= weights[1353];
				12'd1354	: data <= weights[1354];
				12'd1355	: data <= weights[1355];
				12'd1356	: data <= weights[1356];
				12'd1357	: data <= weights[1357];
				12'd1358	: data <= weights[1358];
				12'd1359	: data <= weights[1359];
				12'd1360	: data <= weights[1360];
				12'd1361	: data <= weights[1361];
				12'd1362	: data <= weights[1362];
				12'd1363	: data <= weights[1363];
				12'd1364	: data <= weights[1364];
				12'd1365	: data <= weights[1365];
				12'd1366	: data <= weights[1366];
				12'd1367	: data <= weights[1367];
				12'd1368	: data <= weights[1368];
				12'd1369	: data <= weights[1369];
				12'd1370	: data <= weights[1370];
				12'd1371	: data <= weights[1371];
				12'd1372	: data <= weights[1372];
				12'd1373	: data <= weights[1373];
				12'd1374	: data <= weights[1374];
				12'd1375	: data <= weights[1375];
				12'd1376	: data <= weights[1376];
				12'd1377	: data <= weights[1377];
				12'd1378	: data <= weights[1378];
				12'd1379	: data <= weights[1379];
				12'd1380	: data <= weights[1380];
				12'd1381	: data <= weights[1381];
				12'd1382	: data <= weights[1382];
				12'd1383	: data <= weights[1383];
				12'd1384	: data <= weights[1384];
				12'd1385	: data <= weights[1385];
				12'd1386	: data <= weights[1386];
				12'd1387	: data <= weights[1387];
				12'd1388	: data <= weights[1388];
				12'd1389	: data <= weights[1389];
				12'd1390	: data <= weights[1390];
				12'd1391	: data <= weights[1391];
				12'd1392	: data <= weights[1392];
				12'd1393	: data <= weights[1393];
				12'd1394	: data <= weights[1394];
				12'd1395	: data <= weights[1395];
				12'd1396	: data <= weights[1396];
				12'd1397	: data <= weights[1397];
				12'd1398	: data <= weights[1398];
				12'd1399	: data <= weights[1399];
				12'd1400	: data <= weights[1400];
				12'd1401	: data <= weights[1401];
				12'd1402	: data <= weights[1402];
				12'd1403	: data <= weights[1403];
				12'd1404	: data <= weights[1404];
				12'd1405	: data <= weights[1405];
				12'd1406	: data <= weights[1406];
				12'd1407	: data <= weights[1407];
				12'd1408	: data <= weights[1408];
				12'd1409	: data <= weights[1409];
				12'd1410	: data <= weights[1410];
				12'd1411	: data <= weights[1411];
				12'd1412	: data <= weights[1412];
				12'd1413	: data <= weights[1413];
				12'd1414	: data <= weights[1414];
				12'd1415	: data <= weights[1415];
				12'd1416	: data <= weights[1416];
				12'd1417	: data <= weights[1417];
				12'd1418	: data <= weights[1418];
				12'd1419	: data <= weights[1419];
				12'd1420	: data <= weights[1420];
				12'd1421	: data <= weights[1421];
				12'd1422	: data <= weights[1422];
				12'd1423	: data <= weights[1423];
				12'd1424	: data <= weights[1424];
				12'd1425	: data <= weights[1425];
				12'd1426	: data <= weights[1426];
				12'd1427	: data <= weights[1427];
				12'd1428	: data <= weights[1428];
				12'd1429	: data <= weights[1429];
				12'd1430	: data <= weights[1430];
				12'd1431	: data <= weights[1431];
				12'd1432	: data <= weights[1432];
				12'd1433	: data <= weights[1433];
				12'd1434	: data <= weights[1434];
				12'd1435	: data <= weights[1435];
				12'd1436	: data <= weights[1436];
				12'd1437	: data <= weights[1437];
				12'd1438	: data <= weights[1438];
				12'd1439	: data <= weights[1439];
				12'd1440	: data <= weights[1440];
				12'd1441	: data <= weights[1441];
				12'd1442	: data <= weights[1442];
				12'd1443	: data <= weights[1443];
				12'd1444	: data <= weights[1444];
				12'd1445	: data <= weights[1445];
				12'd1446	: data <= weights[1446];
				12'd1447	: data <= weights[1447];
				12'd1448	: data <= weights[1448];
				12'd1449	: data <= weights[1449];
				12'd1450	: data <= weights[1450];
				12'd1451	: data <= weights[1451];
				12'd1452	: data <= weights[1452];
				12'd1453	: data <= weights[1453];
				12'd1454	: data <= weights[1454];
				12'd1455	: data <= weights[1455];
				12'd1456	: data <= weights[1456];
				12'd1457	: data <= weights[1457];
				12'd1458	: data <= weights[1458];
				12'd1459	: data <= weights[1459];
				12'd1460	: data <= weights[1460];
				12'd1461	: data <= weights[1461];
				12'd1462	: data <= weights[1462];
				12'd1463	: data <= weights[1463];
				12'd1464	: data <= weights[1464];
				12'd1465	: data <= weights[1465];
				12'd1466	: data <= weights[1466];
				12'd1467	: data <= weights[1467];
				12'd1468	: data <= weights[1468];
				12'd1469	: data <= weights[1469];
				12'd1470	: data <= weights[1470];
				12'd1471	: data <= weights[1471];
				12'd1472	: data <= weights[1472];
				12'd1473	: data <= weights[1473];
				12'd1474	: data <= weights[1474];
				12'd1475	: data <= weights[1475];
				12'd1476	: data <= weights[1476];
				12'd1477	: data <= weights[1477];
				12'd1478	: data <= weights[1478];
				12'd1479	: data <= weights[1479];
				12'd1480	: data <= weights[1480];
				12'd1481	: data <= weights[1481];
				12'd1482	: data <= weights[1482];
				12'd1483	: data <= weights[1483];
				12'd1484	: data <= weights[1484];
				12'd1485	: data <= weights[1485];
				12'd1486	: data <= weights[1486];
				12'd1487	: data <= weights[1487];
				12'd1488	: data <= weights[1488];
				12'd1489	: data <= weights[1489];
				12'd1490	: data <= weights[1490];
				12'd1491	: data <= weights[1491];
				12'd1492	: data <= weights[1492];
				12'd1493	: data <= weights[1493];
				12'd1494	: data <= weights[1494];
				12'd1495	: data <= weights[1495];
				12'd1496	: data <= weights[1496];
				12'd1497	: data <= weights[1497];
				12'd1498	: data <= weights[1498];
				12'd1499	: data <= weights[1499];
				12'd1500	: data <= weights[1500];
				12'd1501	: data <= weights[1501];
				12'd1502	: data <= weights[1502];
				12'd1503	: data <= weights[1503];
				12'd1504	: data <= weights[1504];
				12'd1505	: data <= weights[1505];
				12'd1506	: data <= weights[1506];
				12'd1507	: data <= weights[1507];
				12'd1508	: data <= weights[1508];
				12'd1509	: data <= weights[1509];
				12'd1510	: data <= weights[1510];
				12'd1511	: data <= weights[1511];
				12'd1512	: data <= weights[1512];
				12'd1513	: data <= weights[1513];
				12'd1514	: data <= weights[1514];
				12'd1515	: data <= weights[1515];
				12'd1516	: data <= weights[1516];
				12'd1517	: data <= weights[1517];
				12'd1518	: data <= weights[1518];
				12'd1519	: data <= weights[1519];
				12'd1520	: data <= weights[1520];
				12'd1521	: data <= weights[1521];
				12'd1522	: data <= weights[1522];
				12'd1523	: data <= weights[1523];
				12'd1524	: data <= weights[1524];
				12'd1525	: data <= weights[1525];
				12'd1526	: data <= weights[1526];
				12'd1527	: data <= weights[1527];
				12'd1528	: data <= weights[1528];
				12'd1529	: data <= weights[1529];
				12'd1530	: data <= weights[1530];
				12'd1531	: data <= weights[1531];
				12'd1532	: data <= weights[1532];
				12'd1533	: data <= weights[1533];
				12'd1534	: data <= weights[1534];
				12'd1535	: data <= weights[1535];
				12'd1536	: data <= weights[1536];
				12'd1537	: data <= weights[1537];
				12'd1538	: data <= weights[1538];
				12'd1539	: data <= weights[1539];
				12'd1540	: data <= weights[1540];
				12'd1541	: data <= weights[1541];
				12'd1542	: data <= weights[1542];
				12'd1543	: data <= weights[1543];
				12'd1544	: data <= weights[1544];
				12'd1545	: data <= weights[1545];
				12'd1546	: data <= weights[1546];
				12'd1547	: data <= weights[1547];
				12'd1548	: data <= weights[1548];
				12'd1549	: data <= weights[1549];
				12'd1550	: data <= weights[1550];
				12'd1551	: data <= weights[1551];
				12'd1552	: data <= weights[1552];
				12'd1553	: data <= weights[1553];
				12'd1554	: data <= weights[1554];
				12'd1555	: data <= weights[1555];
				12'd1556	: data <= weights[1556];
				12'd1557	: data <= weights[1557];
				12'd1558	: data <= weights[1558];
				12'd1559	: data <= weights[1559];
				12'd1560	: data <= weights[1560];
				12'd1561	: data <= weights[1561];
				12'd1562	: data <= weights[1562];
				12'd1563	: data <= weights[1563];
				12'd1564	: data <= weights[1564];
				12'd1565	: data <= weights[1565];
				12'd1566	: data <= weights[1566];
				12'd1567	: data <= weights[1567];
				12'd1568	: data <= weights[1568];
				12'd1569	: data <= weights[1569];
				12'd1570	: data <= weights[1570];
				12'd1571	: data <= weights[1571];
				12'd1572	: data <= weights[1572];
				12'd1573	: data <= weights[1573];
				12'd1574	: data <= weights[1574];
				12'd1575	: data <= weights[1575];
				12'd1576	: data <= weights[1576];
				12'd1577	: data <= weights[1577];
				12'd1578	: data <= weights[1578];
				12'd1579	: data <= weights[1579];
				12'd1580	: data <= weights[1580];
				12'd1581	: data <= weights[1581];
				12'd1582	: data <= weights[1582];
				12'd1583	: data <= weights[1583];
				12'd1584	: data <= weights[1584];
				12'd1585	: data <= weights[1585];
				12'd1586	: data <= weights[1586];
				12'd1587	: data <= weights[1587];
				12'd1588	: data <= weights[1588];
				12'd1589	: data <= weights[1589];
				12'd1590	: data <= weights[1590];
				12'd1591	: data <= weights[1591];
				12'd1592	: data <= weights[1592];
				12'd1593	: data <= weights[1593];
				12'd1594	: data <= weights[1594];
				12'd1595	: data <= weights[1595];
				12'd1596	: data <= weights[1596];
				12'd1597	: data <= weights[1597];
				12'd1598	: data <= weights[1598];
				12'd1599	: data <= weights[1599];
				12'd1600	: data <= weights[1600];
				12'd1601	: data <= weights[1601];
				12'd1602	: data <= weights[1602];
				12'd1603	: data <= weights[1603];
				12'd1604	: data <= weights[1604];
				12'd1605	: data <= weights[1605];
				12'd1606	: data <= weights[1606];
				12'd1607	: data <= weights[1607];
				12'd1608	: data <= weights[1608];
				12'd1609	: data <= weights[1609];
				12'd1610	: data <= weights[1610];
				12'd1611	: data <= weights[1611];
				12'd1612	: data <= weights[1612];
				12'd1613	: data <= weights[1613];
				12'd1614	: data <= weights[1614];
				12'd1615	: data <= weights[1615];
				12'd1616	: data <= weights[1616];
				12'd1617	: data <= weights[1617];
				12'd1618	: data <= weights[1618];
				12'd1619	: data <= weights[1619];
				12'd1620	: data <= weights[1620];
				12'd1621	: data <= weights[1621];
				12'd1622	: data <= weights[1622];
				12'd1623	: data <= weights[1623];
				12'd1624	: data <= weights[1624];
				12'd1625	: data <= weights[1625];
				12'd1626	: data <= weights[1626];
				12'd1627	: data <= weights[1627];
				12'd1628	: data <= weights[1628];
				12'd1629	: data <= weights[1629];
				12'd1630	: data <= weights[1630];
				12'd1631	: data <= weights[1631];
				12'd1632	: data <= weights[1632];
				12'd1633	: data <= weights[1633];
				12'd1634	: data <= weights[1634];
				12'd1635	: data <= weights[1635];
				12'd1636	: data <= weights[1636];
				12'd1637	: data <= weights[1637];
				12'd1638	: data <= weights[1638];
				12'd1639	: data <= weights[1639];
				12'd1640	: data <= weights[1640];
				12'd1641	: data <= weights[1641];
				12'd1642	: data <= weights[1642];
				12'd1643	: data <= weights[1643];
				12'd1644	: data <= weights[1644];
				12'd1645	: data <= weights[1645];
				12'd1646	: data <= weights[1646];
				12'd1647	: data <= weights[1647];
				12'd1648	: data <= weights[1648];
				12'd1649	: data <= weights[1649];
				12'd1650	: data <= weights[1650];
				12'd1651	: data <= weights[1651];
				12'd1652	: data <= weights[1652];
				12'd1653	: data <= weights[1653];
				12'd1654	: data <= weights[1654];
				12'd1655	: data <= weights[1655];
				12'd1656	: data <= weights[1656];
				12'd1657	: data <= weights[1657];
				12'd1658	: data <= weights[1658];
				12'd1659	: data <= weights[1659];
				12'd1660	: data <= weights[1660];
				12'd1661	: data <= weights[1661];
				12'd1662	: data <= weights[1662];
				12'd1663	: data <= weights[1663];
				12'd1664	: data <= weights[1664];
				12'd1665	: data <= weights[1665];
				12'd1666	: data <= weights[1666];
				12'd1667	: data <= weights[1667];
				12'd1668	: data <= weights[1668];
				12'd1669	: data <= weights[1669];
				12'd1670	: data <= weights[1670];
				12'd1671	: data <= weights[1671];
				12'd1672	: data <= weights[1672];
				12'd1673	: data <= weights[1673];
				12'd1674	: data <= weights[1674];
				12'd1675	: data <= weights[1675];
				12'd1676	: data <= weights[1676];
				12'd1677	: data <= weights[1677];
				12'd1678	: data <= weights[1678];
				12'd1679	: data <= weights[1679];
				12'd1680	: data <= weights[1680];
				12'd1681	: data <= weights[1681];
				12'd1682	: data <= weights[1682];
				12'd1683	: data <= weights[1683];
				12'd1684	: data <= weights[1684];
				12'd1685	: data <= weights[1685];
				12'd1686	: data <= weights[1686];
				12'd1687	: data <= weights[1687];
				12'd1688	: data <= weights[1688];
				12'd1689	: data <= weights[1689];
				12'd1690	: data <= weights[1690];
				12'd1691	: data <= weights[1691];
				12'd1692	: data <= weights[1692];
				12'd1693	: data <= weights[1693];
				12'd1694	: data <= weights[1694];
				12'd1695	: data <= weights[1695];
				12'd1696	: data <= weights[1696];
				12'd1697	: data <= weights[1697];
				12'd1698	: data <= weights[1698];
				12'd1699	: data <= weights[1699];
				12'd1700	: data <= weights[1700];
				12'd1701	: data <= weights[1701];
				12'd1702	: data <= weights[1702];
				12'd1703	: data <= weights[1703];
				12'd1704	: data <= weights[1704];
				12'd1705	: data <= weights[1705];
				12'd1706	: data <= weights[1706];
				12'd1707	: data <= weights[1707];
				12'd1708	: data <= weights[1708];
				12'd1709	: data <= weights[1709];
				12'd1710	: data <= weights[1710];
				12'd1711	: data <= weights[1711];
				12'd1712	: data <= weights[1712];
				12'd1713	: data <= weights[1713];
				12'd1714	: data <= weights[1714];
				12'd1715	: data <= weights[1715];
				12'd1716	: data <= weights[1716];
				12'd1717	: data <= weights[1717];
				12'd1718	: data <= weights[1718];
				12'd1719	: data <= weights[1719];
				12'd1720	: data <= weights[1720];
				12'd1721	: data <= weights[1721];
				12'd1722	: data <= weights[1722];
				12'd1723	: data <= weights[1723];
				12'd1724	: data <= weights[1724];
				12'd1725	: data <= weights[1725];
				12'd1726	: data <= weights[1726];
				12'd1727	: data <= weights[1727];
				12'd1728	: data <= weights[1728];
				12'd1729	: data <= weights[1729];
				12'd1730	: data <= weights[1730];
				12'd1731	: data <= weights[1731];
				12'd1732	: data <= weights[1732];
				12'd1733	: data <= weights[1733];
				12'd1734	: data <= weights[1734];
				12'd1735	: data <= weights[1735];
				12'd1736	: data <= weights[1736];
				12'd1737	: data <= weights[1737];
				12'd1738	: data <= weights[1738];
				12'd1739	: data <= weights[1739];
				12'd1740	: data <= weights[1740];
				12'd1741	: data <= weights[1741];
				12'd1742	: data <= weights[1742];
				12'd1743	: data <= weights[1743];
				12'd1744	: data <= weights[1744];
				12'd1745	: data <= weights[1745];
				12'd1746	: data <= weights[1746];
				12'd1747	: data <= weights[1747];
				12'd1748	: data <= weights[1748];
				12'd1749	: data <= weights[1749];
				12'd1750	: data <= weights[1750];
				12'd1751	: data <= weights[1751];
				12'd1752	: data <= weights[1752];
				12'd1753	: data <= weights[1753];
				12'd1754	: data <= weights[1754];
				12'd1755	: data <= weights[1755];
				12'd1756	: data <= weights[1756];
				12'd1757	: data <= weights[1757];
				12'd1758	: data <= weights[1758];
				12'd1759	: data <= weights[1759];
				12'd1760	: data <= weights[1760];
				12'd1761	: data <= weights[1761];
				12'd1762	: data <= weights[1762];
				12'd1763	: data <= weights[1763];
				12'd1764	: data <= weights[1764];
				12'd1765	: data <= weights[1765];
				12'd1766	: data <= weights[1766];
				12'd1767	: data <= weights[1767];
				12'd1768	: data <= weights[1768];
				12'd1769	: data <= weights[1769];
				12'd1770	: data <= weights[1770];
				12'd1771	: data <= weights[1771];
				12'd1772	: data <= weights[1772];
				12'd1773	: data <= weights[1773];
				12'd1774	: data <= weights[1774];
				12'd1775	: data <= weights[1775];
				12'd1776	: data <= weights[1776];
				12'd1777	: data <= weights[1777];
				12'd1778	: data <= weights[1778];
				12'd1779	: data <= weights[1779];
				12'd1780	: data <= weights[1780];
				12'd1781	: data <= weights[1781];
				12'd1782	: data <= weights[1782];
				12'd1783	: data <= weights[1783];
				12'd1784	: data <= weights[1784];
				12'd1785	: data <= weights[1785];
				12'd1786	: data <= weights[1786];
				12'd1787	: data <= weights[1787];
				12'd1788	: data <= weights[1788];
				12'd1789	: data <= weights[1789];
				12'd1790	: data <= weights[1790];
				12'd1791	: data <= weights[1791];
				12'd1792	: data <= weights[1792];
				12'd1793	: data <= weights[1793];
				12'd1794	: data <= weights[1794];
				12'd1795	: data <= weights[1795];
				12'd1796	: data <= weights[1796];
				12'd1797	: data <= weights[1797];
				12'd1798	: data <= weights[1798];
				12'd1799	: data <= weights[1799];
				12'd1800	: data <= weights[1800];
				12'd1801	: data <= weights[1801];
				12'd1802	: data <= weights[1802];
				12'd1803	: data <= weights[1803];
				12'd1804	: data <= weights[1804];
				12'd1805	: data <= weights[1805];
				12'd1806	: data <= weights[1806];
				12'd1807	: data <= weights[1807];
				12'd1808	: data <= weights[1808];
				12'd1809	: data <= weights[1809];
				12'd1810	: data <= weights[1810];
				12'd1811	: data <= weights[1811];
				12'd1812	: data <= weights[1812];
				12'd1813	: data <= weights[1813];
				12'd1814	: data <= weights[1814];
				12'd1815	: data <= weights[1815];
				12'd1816	: data <= weights[1816];
				12'd1817	: data <= weights[1817];
				12'd1818	: data <= weights[1818];
				12'd1819	: data <= weights[1819];
				12'd1820	: data <= weights[1820];
				12'd1821	: data <= weights[1821];
				12'd1822	: data <= weights[1822];
				12'd1823	: data <= weights[1823];
				12'd1824	: data <= weights[1824];
				12'd1825	: data <= weights[1825];
				12'd1826	: data <= weights[1826];
				12'd1827	: data <= weights[1827];
				12'd1828	: data <= weights[1828];
				12'd1829	: data <= weights[1829];
				12'd1830	: data <= weights[1830];
				12'd1831	: data <= weights[1831];
				12'd1832	: data <= weights[1832];
				12'd1833	: data <= weights[1833];
				12'd1834	: data <= weights[1834];
				12'd1835	: data <= weights[1835];
				12'd1836	: data <= weights[1836];
				12'd1837	: data <= weights[1837];
				12'd1838	: data <= weights[1838];
				12'd1839	: data <= weights[1839];
				12'd1840	: data <= weights[1840];
				12'd1841	: data <= weights[1841];
				12'd1842	: data <= weights[1842];
				12'd1843	: data <= weights[1843];
				12'd1844	: data <= weights[1844];
				12'd1845	: data <= weights[1845];
				12'd1846	: data <= weights[1846];
				12'd1847	: data <= weights[1847];
				12'd1848	: data <= weights[1848];
				12'd1849	: data <= weights[1849];
				12'd1850	: data <= weights[1850];
				12'd1851	: data <= weights[1851];
				12'd1852	: data <= weights[1852];
				12'd1853	: data <= weights[1853];
				12'd1854	: data <= weights[1854];
				12'd1855	: data <= weights[1855];
				12'd1856	: data <= weights[1856];
				12'd1857	: data <= weights[1857];
				12'd1858	: data <= weights[1858];
				12'd1859	: data <= weights[1859];
				12'd1860	: data <= weights[1860];
				12'd1861	: data <= weights[1861];
				12'd1862	: data <= weights[1862];
				12'd1863	: data <= weights[1863];
				12'd1864	: data <= weights[1864];
				12'd1865	: data <= weights[1865];
				12'd1866	: data <= weights[1866];
				12'd1867	: data <= weights[1867];
				12'd1868	: data <= weights[1868];
				12'd1869	: data <= weights[1869];
				12'd1870	: data <= weights[1870];
				12'd1871	: data <= weights[1871];
				12'd1872	: data <= weights[1872];
				12'd1873	: data <= weights[1873];
				12'd1874	: data <= weights[1874];
				12'd1875	: data <= weights[1875];
				12'd1876	: data <= weights[1876];
				12'd1877	: data <= weights[1877];
				12'd1878	: data <= weights[1878];
				12'd1879	: data <= weights[1879];
				12'd1880	: data <= weights[1880];
				12'd1881	: data <= weights[1881];
				12'd1882	: data <= weights[1882];
				12'd1883	: data <= weights[1883];
				12'd1884	: data <= weights[1884];
				12'd1885	: data <= weights[1885];
				12'd1886	: data <= weights[1886];
				12'd1887	: data <= weights[1887];
				12'd1888	: data <= weights[1888];
				12'd1889	: data <= weights[1889];
				12'd1890	: data <= weights[1890];
				12'd1891	: data <= weights[1891];
				12'd1892	: data <= weights[1892];
				12'd1893	: data <= weights[1893];
				12'd1894	: data <= weights[1894];
				12'd1895	: data <= weights[1895];
				12'd1896	: data <= weights[1896];
				12'd1897	: data <= weights[1897];
				12'd1898	: data <= weights[1898];
				12'd1899	: data <= weights[1899];
				12'd1900	: data <= weights[1900];
				12'd1901	: data <= weights[1901];
				12'd1902	: data <= weights[1902];
				12'd1903	: data <= weights[1903];
				12'd1904	: data <= weights[1904];
				12'd1905	: data <= weights[1905];
				12'd1906	: data <= weights[1906];
				12'd1907	: data <= weights[1907];
				12'd1908	: data <= weights[1908];
				12'd1909	: data <= weights[1909];
				12'd1910	: data <= weights[1910];
				12'd1911	: data <= weights[1911];
				12'd1912	: data <= weights[1912];
				12'd1913	: data <= weights[1913];
				12'd1914	: data <= weights[1914];
				12'd1915	: data <= weights[1915];
				12'd1916	: data <= weights[1916];
				12'd1917	: data <= weights[1917];
				12'd1918	: data <= weights[1918];
				12'd1919	: data <= weights[1919];
				12'd1920	: data <= weights[1920];
				12'd1921	: data <= weights[1921];
				12'd1922	: data <= weights[1922];
				12'd1923	: data <= weights[1923];
				12'd1924	: data <= weights[1924];
				12'd1925	: data <= weights[1925];
				12'd1926	: data <= weights[1926];
				12'd1927	: data <= weights[1927];
				12'd1928	: data <= weights[1928];
				12'd1929	: data <= weights[1929];
				12'd1930	: data <= weights[1930];
				12'd1931	: data <= weights[1931];
				12'd1932	: data <= weights[1932];
				12'd1933	: data <= weights[1933];
				12'd1934	: data <= weights[1934];
				12'd1935	: data <= weights[1935];
				12'd1936	: data <= weights[1936];
				12'd1937	: data <= weights[1937];
				12'd1938	: data <= weights[1938];
				12'd1939	: data <= weights[1939];
				12'd1940	: data <= weights[1940];
				12'd1941	: data <= weights[1941];
				12'd1942	: data <= weights[1942];
				12'd1943	: data <= weights[1943];
				12'd1944	: data <= weights[1944];
				12'd1945	: data <= weights[1945];
				12'd1946	: data <= weights[1946];
				12'd1947	: data <= weights[1947];
				12'd1948	: data <= weights[1948];
				12'd1949	: data <= weights[1949];
				12'd1950	: data <= weights[1950];
				12'd1951	: data <= weights[1951];
				12'd1952	: data <= weights[1952];
				12'd1953	: data <= weights[1953];
				12'd1954	: data <= weights[1954];
				12'd1955	: data <= weights[1955];
				12'd1956	: data <= weights[1956];
				12'd1957	: data <= weights[1957];
				12'd1958	: data <= weights[1958];
				12'd1959	: data <= weights[1959];
				12'd1960	: data <= weights[1960];
				12'd1961	: data <= weights[1961];
				12'd1962	: data <= weights[1962];
				12'd1963	: data <= weights[1963];
				12'd1964	: data <= weights[1964];
				12'd1965	: data <= weights[1965];
				12'd1966	: data <= weights[1966];
				12'd1967	: data <= weights[1967];
				12'd1968	: data <= weights[1968];
				12'd1969	: data <= weights[1969];
				12'd1970	: data <= weights[1970];
				12'd1971	: data <= weights[1971];
				12'd1972	: data <= weights[1972];
				12'd1973	: data <= weights[1973];
				12'd1974	: data <= weights[1974];
				12'd1975	: data <= weights[1975];
				12'd1976	: data <= weights[1976];
				12'd1977	: data <= weights[1977];
				12'd1978	: data <= weights[1978];
				12'd1979	: data <= weights[1979];
				12'd1980	: data <= weights[1980];
				12'd1981	: data <= weights[1981];
				12'd1982	: data <= weights[1982];
				12'd1983	: data <= weights[1983];
				12'd1984	: data <= weights[1984];
				12'd1985	: data <= weights[1985];
				12'd1986	: data <= weights[1986];
				12'd1987	: data <= weights[1987];
				12'd1988	: data <= weights[1988];
				12'd1989	: data <= weights[1989];
				12'd1990	: data <= weights[1990];
				12'd1991	: data <= weights[1991];
				12'd1992	: data <= weights[1992];
				12'd1993	: data <= weights[1993];
				12'd1994	: data <= weights[1994];
				12'd1995	: data <= weights[1995];
				12'd1996	: data <= weights[1996];
				12'd1997	: data <= weights[1997];
				12'd1998	: data <= weights[1998];
				12'd1999	: data <= weights[1999];
				12'd2000	: data <= weights[2000];
				12'd2001	: data <= weights[2001];
				12'd2002	: data <= weights[2002];
				12'd2003	: data <= weights[2003];
				12'd2004	: data <= weights[2004];
				12'd2005	: data <= weights[2005];
				12'd2006	: data <= weights[2006];
				12'd2007	: data <= weights[2007];
				12'd2008	: data <= weights[2008];
				12'd2009	: data <= weights[2009];
				12'd2010	: data <= weights[2010];
				12'd2011	: data <= weights[2011];
				12'd2012	: data <= weights[2012];
				12'd2013	: data <= weights[2013];
				12'd2014	: data <= weights[2014];
				12'd2015	: data <= weights[2015];
				12'd2016	: data <= weights[2016];
				12'd2017	: data <= weights[2017];
				12'd2018	: data <= weights[2018];
				12'd2019	: data <= weights[2019];
				12'd2020	: data <= weights[2020];
				12'd2021	: data <= weights[2021];
				12'd2022	: data <= weights[2022];
				12'd2023	: data <= weights[2023];
				12'd2024	: data <= weights[2024];
				12'd2025	: data <= weights[2025];
				12'd2026	: data <= weights[2026];
				12'd2027	: data <= weights[2027];
				12'd2028	: data <= weights[2028];
				12'd2029	: data <= weights[2029];
				12'd2030	: data <= weights[2030];
				12'd2031	: data <= weights[2031];
				12'd2032	: data <= weights[2032];
				12'd2033	: data <= weights[2033];
				12'd2034	: data <= weights[2034];
				12'd2035	: data <= weights[2035];
				12'd2036	: data <= weights[2036];
				12'd2037	: data <= weights[2037];
				12'd2038	: data <= weights[2038];
				12'd2039	: data <= weights[2039];
				12'd2040	: data <= weights[2040];
				12'd2041	: data <= weights[2041];
				12'd2042	: data <= weights[2042];
				12'd2043	: data <= weights[2043];
				12'd2044	: data <= weights[2044];
				12'd2045	: data <= weights[2045];
				12'd2046	: data <= weights[2046];
				12'd2047	: data <= weights[2047];
				12'd2048	: data <= weights[2048];
				12'd2049	: data <= weights[2049];
				12'd2050	: data <= weights[2050];
				12'd2051	: data <= weights[2051];
				12'd2052	: data <= weights[2052];
				12'd2053	: data <= weights[2053];
				12'd2054	: data <= weights[2054];
				12'd2055	: data <= weights[2055];
				12'd2056	: data <= weights[2056];
				12'd2057	: data <= weights[2057];
				12'd2058	: data <= weights[2058];
				12'd2059	: data <= weights[2059];
				12'd2060	: data <= weights[2060];
				12'd2061	: data <= weights[2061];
				12'd2062	: data <= weights[2062];
				12'd2063	: data <= weights[2063];
				12'd2064	: data <= weights[2064];
				12'd2065	: data <= weights[2065];
				12'd2066	: data <= weights[2066];
				12'd2067	: data <= weights[2067];
				12'd2068	: data <= weights[2068];
				12'd2069	: data <= weights[2069];
				12'd2070	: data <= weights[2070];
				12'd2071	: data <= weights[2071];
				12'd2072	: data <= weights[2072];
				12'd2073	: data <= weights[2073];
				12'd2074	: data <= weights[2074];
				12'd2075	: data <= weights[2075];
				12'd2076	: data <= weights[2076];
				12'd2077	: data <= weights[2077];
				12'd2078	: data <= weights[2078];
				12'd2079	: data <= weights[2079];
				12'd2080	: data <= weights[2080];
				12'd2081	: data <= weights[2081];
				12'd2082	: data <= weights[2082];
				12'd2083	: data <= weights[2083];
				12'd2084	: data <= weights[2084];
				12'd2085	: data <= weights[2085];
				12'd2086	: data <= weights[2086];
				12'd2087	: data <= weights[2087];
				12'd2088	: data <= weights[2088];
				12'd2089	: data <= weights[2089];
				12'd2090	: data <= weights[2090];
				12'd2091	: data <= weights[2091];
				12'd2092	: data <= weights[2092];
				12'd2093	: data <= weights[2093];
				12'd2094	: data <= weights[2094];
				12'd2095	: data <= weights[2095];
				12'd2096	: data <= weights[2096];
				12'd2097	: data <= weights[2097];
				12'd2098	: data <= weights[2098];
				12'd2099	: data <= weights[2099];
				12'd2100	: data <= weights[2100];
				12'd2101	: data <= weights[2101];
				12'd2102	: data <= weights[2102];
				12'd2103	: data <= weights[2103];
				12'd2104	: data <= weights[2104];
				12'd2105	: data <= weights[2105];
				12'd2106	: data <= weights[2106];
				12'd2107	: data <= weights[2107];
				12'd2108	: data <= weights[2108];
				12'd2109	: data <= weights[2109];
				12'd2110	: data <= weights[2110];
				12'd2111	: data <= weights[2111];
				12'd2112	: data <= weights[2112];
				12'd2113	: data <= weights[2113];
				12'd2114	: data <= weights[2114];
				12'd2115	: data <= weights[2115];
				12'd2116	: data <= weights[2116];
				12'd2117	: data <= weights[2117];
				12'd2118	: data <= weights[2118];
				12'd2119	: data <= weights[2119];
				12'd2120	: data <= weights[2120];
				12'd2121	: data <= weights[2121];
				12'd2122	: data <= weights[2122];
				12'd2123	: data <= weights[2123];
				12'd2124	: data <= weights[2124];
				12'd2125	: data <= weights[2125];
				12'd2126	: data <= weights[2126];
				12'd2127	: data <= weights[2127];
				12'd2128	: data <= weights[2128];
				12'd2129	: data <= weights[2129];
				12'd2130	: data <= weights[2130];
				12'd2131	: data <= weights[2131];
				12'd2132	: data <= weights[2132];
				12'd2133	: data <= weights[2133];
				12'd2134	: data <= weights[2134];
				12'd2135	: data <= weights[2135];
				12'd2136	: data <= weights[2136];
				12'd2137	: data <= weights[2137];
				12'd2138	: data <= weights[2138];
				12'd2139	: data <= weights[2139];
				12'd2140	: data <= weights[2140];
				12'd2141	: data <= weights[2141];
				12'd2142	: data <= weights[2142];
				12'd2143	: data <= weights[2143];
				12'd2144	: data <= weights[2144];
				12'd2145	: data <= weights[2145];
				12'd2146	: data <= weights[2146];
				12'd2147	: data <= weights[2147];
				12'd2148	: data <= weights[2148];
				12'd2149	: data <= weights[2149];
				12'd2150	: data <= weights[2150];
				12'd2151	: data <= weights[2151];
				12'd2152	: data <= weights[2152];
				12'd2153	: data <= weights[2153];
				12'd2154	: data <= weights[2154];
				12'd2155	: data <= weights[2155];
				12'd2156	: data <= weights[2156];
				12'd2157	: data <= weights[2157];
				12'd2158	: data <= weights[2158];
				12'd2159	: data <= weights[2159];
				12'd2160	: data <= weights[2160];
				12'd2161	: data <= weights[2161];
				12'd2162	: data <= weights[2162];
				12'd2163	: data <= weights[2163];
				12'd2164	: data <= weights[2164];
				12'd2165	: data <= weights[2165];
				12'd2166	: data <= weights[2166];
				12'd2167	: data <= weights[2167];
				12'd2168	: data <= weights[2168];
				12'd2169	: data <= weights[2169];
				12'd2170	: data <= weights[2170];
				12'd2171	: data <= weights[2171];
				12'd2172	: data <= weights[2172];
				12'd2173	: data <= weights[2173];
				12'd2174	: data <= weights[2174];
				12'd2175	: data <= weights[2175];
				12'd2176	: data <= weights[2176];
				12'd2177	: data <= weights[2177];
				12'd2178	: data <= weights[2178];
				12'd2179	: data <= weights[2179];
				12'd2180	: data <= weights[2180];
				12'd2181	: data <= weights[2181];
				12'd2182	: data <= weights[2182];
				12'd2183	: data <= weights[2183];
				12'd2184	: data <= weights[2184];
				12'd2185	: data <= weights[2185];
				12'd2186	: data <= weights[2186];
				12'd2187	: data <= weights[2187];
				12'd2188	: data <= weights[2188];
				12'd2189	: data <= weights[2189];
				12'd2190	: data <= weights[2190];
				12'd2191	: data <= weights[2191];
				12'd2192	: data <= weights[2192];
				12'd2193	: data <= weights[2193];
				12'd2194	: data <= weights[2194];
				12'd2195	: data <= weights[2195];
				12'd2196	: data <= weights[2196];
				12'd2197	: data <= weights[2197];
				12'd2198	: data <= weights[2198];
				12'd2199	: data <= weights[2199];
				12'd2200	: data <= weights[2200];
				12'd2201	: data <= weights[2201];
				12'd2202	: data <= weights[2202];
				12'd2203	: data <= weights[2203];
				12'd2204	: data <= weights[2204];
				12'd2205	: data <= weights[2205];
				12'd2206	: data <= weights[2206];
				12'd2207	: data <= weights[2207];
				12'd2208	: data <= weights[2208];
				12'd2209	: data <= weights[2209];
				12'd2210	: data <= weights[2210];
				12'd2211	: data <= weights[2211];
				12'd2212	: data <= weights[2212];
				12'd2213	: data <= weights[2213];
				12'd2214	: data <= weights[2214];
				12'd2215	: data <= weights[2215];
				12'd2216	: data <= weights[2216];
				12'd2217	: data <= weights[2217];
				12'd2218	: data <= weights[2218];
				12'd2219	: data <= weights[2219];
				12'd2220	: data <= weights[2220];
				12'd2221	: data <= weights[2221];
				12'd2222	: data <= weights[2222];
				12'd2223	: data <= weights[2223];
				12'd2224	: data <= weights[2224];
				12'd2225	: data <= weights[2225];
				12'd2226	: data <= weights[2226];
				12'd2227	: data <= weights[2227];
				12'd2228	: data <= weights[2228];
				12'd2229	: data <= weights[2229];
				12'd2230	: data <= weights[2230];
				12'd2231	: data <= weights[2231];
				12'd2232	: data <= weights[2232];
				12'd2233	: data <= weights[2233];
				12'd2234	: data <= weights[2234];
				12'd2235	: data <= weights[2235];
				12'd2236	: data <= weights[2236];
				12'd2237	: data <= weights[2237];
				12'd2238	: data <= weights[2238];
				12'd2239	: data <= weights[2239];
				12'd2240	: data <= weights[2240];
				12'd2241	: data <= weights[2241];
				12'd2242	: data <= weights[2242];
				12'd2243	: data <= weights[2243];
				12'd2244	: data <= weights[2244];
				12'd2245	: data <= weights[2245];
				12'd2246	: data <= weights[2246];
				12'd2247	: data <= weights[2247];
				12'd2248	: data <= weights[2248];
				12'd2249	: data <= weights[2249];
				12'd2250	: data <= weights[2250];
				12'd2251	: data <= weights[2251];
				12'd2252	: data <= weights[2252];
				12'd2253	: data <= weights[2253];
				12'd2254	: data <= weights[2254];
				12'd2255	: data <= weights[2255];
				12'd2256	: data <= weights[2256];
				12'd2257	: data <= weights[2257];
				12'd2258	: data <= weights[2258];
				12'd2259	: data <= weights[2259];
				12'd2260	: data <= weights[2260];
				12'd2261	: data <= weights[2261];
				12'd2262	: data <= weights[2262];
				12'd2263	: data <= weights[2263];
				12'd2264	: data <= weights[2264];
				12'd2265	: data <= weights[2265];
				12'd2266	: data <= weights[2266];
				12'd2267	: data <= weights[2267];
				12'd2268	: data <= weights[2268];
				12'd2269	: data <= weights[2269];
				12'd2270	: data <= weights[2270];
				12'd2271	: data <= weights[2271];
				12'd2272	: data <= weights[2272];
				12'd2273	: data <= weights[2273];
				12'd2274	: data <= weights[2274];
				12'd2275	: data <= weights[2275];
				12'd2276	: data <= weights[2276];
				12'd2277	: data <= weights[2277];
				12'd2278	: data <= weights[2278];
				12'd2279	: data <= weights[2279];
				12'd2280	: data <= weights[2280];
				12'd2281	: data <= weights[2281];
				12'd2282	: data <= weights[2282];
				12'd2283	: data <= weights[2283];
				12'd2284	: data <= weights[2284];
				12'd2285	: data <= weights[2285];
				12'd2286	: data <= weights[2286];
				12'd2287	: data <= weights[2287];
				12'd2288	: data <= weights[2288];
				12'd2289	: data <= weights[2289];
				12'd2290	: data <= weights[2290];
				12'd2291	: data <= weights[2291];
				12'd2292	: data <= weights[2292];
				12'd2293	: data <= weights[2293];
				12'd2294	: data <= weights[2294];
				12'd2295	: data <= weights[2295];
				12'd2296	: data <= weights[2296];
				12'd2297	: data <= weights[2297];
				12'd2298	: data <= weights[2298];
				12'd2299	: data <= weights[2299];
				12'd2300	: data <= weights[2300];
				12'd2301	: data <= weights[2301];
				12'd2302	: data <= weights[2302];
				12'd2303	: data <= weights[2303];
				12'd2304	: data <= weights[2304];
				12'd2305	: data <= weights[2305];
				12'd2306	: data <= weights[2306];
				12'd2307	: data <= weights[2307];
				12'd2308	: data <= weights[2308];
				12'd2309	: data <= weights[2309];
				12'd2310	: data <= weights[2310];
				12'd2311	: data <= weights[2311];
				12'd2312	: data <= weights[2312];
				12'd2313	: data <= weights[2313];
				12'd2314	: data <= weights[2314];
				12'd2315	: data <= weights[2315];
				12'd2316	: data <= weights[2316];
				12'd2317	: data <= weights[2317];
				12'd2318	: data <= weights[2318];
				12'd2319	: data <= weights[2319];
				12'd2320	: data <= weights[2320];
				12'd2321	: data <= weights[2321];
				12'd2322	: data <= weights[2322];
				12'd2323	: data <= weights[2323];
				12'd2324	: data <= weights[2324];
				12'd2325	: data <= weights[2325];
				12'd2326	: data <= weights[2326];
				12'd2327	: data <= weights[2327];
				12'd2328	: data <= weights[2328];
				12'd2329	: data <= weights[2329];
				12'd2330	: data <= weights[2330];
				12'd2331	: data <= weights[2331];
				12'd2332	: data <= weights[2332];
				12'd2333	: data <= weights[2333];
				12'd2334	: data <= weights[2334];
				12'd2335	: data <= weights[2335];
				12'd2336	: data <= weights[2336];
				12'd2337	: data <= weights[2337];
				12'd2338	: data <= weights[2338];
				12'd2339	: data <= weights[2339];
				12'd2340	: data <= weights[2340];
				12'd2341	: data <= weights[2341];
				12'd2342	: data <= weights[2342];
				12'd2343	: data <= weights[2343];
				12'd2344	: data <= weights[2344];
				12'd2345	: data <= weights[2345];
				12'd2346	: data <= weights[2346];
				12'd2347	: data <= weights[2347];
				12'd2348	: data <= weights[2348];
				12'd2349	: data <= weights[2349];
				12'd2350	: data <= weights[2350];
				12'd2351	: data <= weights[2351];
				12'd2352	: data <= weights[2352];
				12'd2353	: data <= weights[2353];
				12'd2354	: data <= weights[2354];
				12'd2355	: data <= weights[2355];
				12'd2356	: data <= weights[2356];
				12'd2357	: data <= weights[2357];
				12'd2358	: data <= weights[2358];
				12'd2359	: data <= weights[2359];
				12'd2360	: data <= weights[2360];
				12'd2361	: data <= weights[2361];
				12'd2362	: data <= weights[2362];
				12'd2363	: data <= weights[2363];
				12'd2364	: data <= weights[2364];
				12'd2365	: data <= weights[2365];
				12'd2366	: data <= weights[2366];
				12'd2367	: data <= weights[2367];
				12'd2368	: data <= weights[2368];
				12'd2369	: data <= weights[2369];
				12'd2370	: data <= weights[2370];
				12'd2371	: data <= weights[2371];
				12'd2372	: data <= weights[2372];
				12'd2373	: data <= weights[2373];
				12'd2374	: data <= weights[2374];
				12'd2375	: data <= weights[2375];
				12'd2376	: data <= weights[2376];
				12'd2377	: data <= weights[2377];
				12'd2378	: data <= weights[2378];
				12'd2379	: data <= weights[2379];
				12'd2380	: data <= weights[2380];
				12'd2381	: data <= weights[2381];
				12'd2382	: data <= weights[2382];
				12'd2383	: data <= weights[2383];
				12'd2384	: data <= weights[2384];
				12'd2385	: data <= weights[2385];
				12'd2386	: data <= weights[2386];
				12'd2387	: data <= weights[2387];
				12'd2388	: data <= weights[2388];
				12'd2389	: data <= weights[2389];
				12'd2390	: data <= weights[2390];
				12'd2391	: data <= weights[2391];
				12'd2392	: data <= weights[2392];
				12'd2393	: data <= weights[2393];
				12'd2394	: data <= weights[2394];
				12'd2395	: data <= weights[2395];
				12'd2396	: data <= weights[2396];
				12'd2397	: data <= weights[2397];
				12'd2398	: data <= weights[2398];
				12'd2399	: data <= weights[2399];
				12'd2400	: data <= weights[2400];
				12'd2401	: data <= weights[2401];
				12'd2402	: data <= weights[2402];
				12'd2403	: data <= weights[2403];
				12'd2404	: data <= weights[2404];
				12'd2405	: data <= weights[2405];
				12'd2406	: data <= weights[2406];
				12'd2407	: data <= weights[2407];
				12'd2408	: data <= weights[2408];
				12'd2409	: data <= weights[2409];
				12'd2410	: data <= weights[2410];
				12'd2411	: data <= weights[2411];
				12'd2412	: data <= weights[2412];
				12'd2413	: data <= weights[2413];
				12'd2414	: data <= weights[2414];
				12'd2415	: data <= weights[2415];
				12'd2416	: data <= weights[2416];
				12'd2417	: data <= weights[2417];
				12'd2418	: data <= weights[2418];
				12'd2419	: data <= weights[2419];
				12'd2420	: data <= weights[2420];
				12'd2421	: data <= weights[2421];
				12'd2422	: data <= weights[2422];
				12'd2423	: data <= weights[2423];
				12'd2424	: data <= weights[2424];
				12'd2425	: data <= weights[2425];
				12'd2426	: data <= weights[2426];
				12'd2427	: data <= weights[2427];
				12'd2428	: data <= weights[2428];
				12'd2429	: data <= weights[2429];
				12'd2430	: data <= weights[2430];
				12'd2431	: data <= weights[2431];
				12'd2432	: data <= weights[2432];
				12'd2433	: data <= weights[2433];
				12'd2434	: data <= weights[2434];
				12'd2435	: data <= weights[2435];
				12'd2436	: data <= weights[2436];
				12'd2437	: data <= weights[2437];
				12'd2438	: data <= weights[2438];
				12'd2439	: data <= weights[2439];
				12'd2440	: data <= weights[2440];
				12'd2441	: data <= weights[2441];
				12'd2442	: data <= weights[2442];
				12'd2443	: data <= weights[2443];
				12'd2444	: data <= weights[2444];
				12'd2445	: data <= weights[2445];
				12'd2446	: data <= weights[2446];
				12'd2447	: data <= weights[2447];
				12'd2448	: data <= weights[2448];
				12'd2449	: data <= weights[2449];
				12'd2450	: data <= weights[2450];
				12'd2451	: data <= weights[2451];
				12'd2452	: data <= weights[2452];
				12'd2453	: data <= weights[2453];
				12'd2454	: data <= weights[2454];
				12'd2455	: data <= weights[2455];
				12'd2456	: data <= weights[2456];
				12'd2457	: data <= weights[2457];
				12'd2458	: data <= weights[2458];
				12'd2459	: data <= weights[2459];
				12'd2460	: data <= weights[2460];
				12'd2461	: data <= weights[2461];
				12'd2462	: data <= weights[2462];
				12'd2463	: data <= weights[2463];
				12'd2464	: data <= weights[2464];
				12'd2465	: data <= weights[2465];
				12'd2466	: data <= weights[2466];
				12'd2467	: data <= weights[2467];
				12'd2468	: data <= weights[2468];
				12'd2469	: data <= weights[2469];
				12'd2470	: data <= weights[2470];
				12'd2471	: data <= weights[2471];
				12'd2472	: data <= weights[2472];
				12'd2473	: data <= weights[2473];
				12'd2474	: data <= weights[2474];
				12'd2475	: data <= weights[2475];
				12'd2476	: data <= weights[2476];
				12'd2477	: data <= weights[2477];
				12'd2478	: data <= weights[2478];
				12'd2479	: data <= weights[2479];
				12'd2480	: data <= weights[2480];
				12'd2481	: data <= weights[2481];
				12'd2482	: data <= weights[2482];
				12'd2483	: data <= weights[2483];
				12'd2484	: data <= weights[2484];
				12'd2485	: data <= weights[2485];
				12'd2486	: data <= weights[2486];
				12'd2487	: data <= weights[2487];
				12'd2488	: data <= weights[2488];
				12'd2489	: data <= weights[2489];
				12'd2490	: data <= weights[2490];
				12'd2491	: data <= weights[2491];
				12'd2492	: data <= weights[2492];
				12'd2493	: data <= weights[2493];
				12'd2494	: data <= weights[2494];
				12'd2495	: data <= weights[2495];
				12'd2496	: data <= weights[2496];
				12'd2497	: data <= weights[2497];
				12'd2498	: data <= weights[2498];
				12'd2499	: data <= weights[2499];
				12'd2500	: data <= weights[2500];
				12'd2501	: data <= weights[2501];
				12'd2502	: data <= weights[2502];
				12'd2503	: data <= weights[2503];
				12'd2504	: data <= weights[2504];
				12'd2505	: data <= weights[2505];
				12'd2506	: data <= weights[2506];
				12'd2507	: data <= weights[2507];
				12'd2508	: data <= weights[2508];
				12'd2509	: data <= weights[2509];
				12'd2510	: data <= weights[2510];
				12'd2511	: data <= weights[2511];
				12'd2512	: data <= weights[2512];
				12'd2513	: data <= weights[2513];
				12'd2514	: data <= weights[2514];
				12'd2515	: data <= weights[2515];
				12'd2516	: data <= weights[2516];
				12'd2517	: data <= weights[2517];
				12'd2518	: data <= weights[2518];
				12'd2519	: data <= weights[2519];
				12'd2520	: data <= weights[2520];
				12'd2521	: data <= weights[2521];
				12'd2522	: data <= weights[2522];
				12'd2523	: data <= weights[2523];
				12'd2524	: data <= weights[2524];
				12'd2525	: data <= weights[2525];
				12'd2526	: data <= weights[2526];
				12'd2527	: data <= weights[2527];
				12'd2528	: data <= weights[2528];
				12'd2529	: data <= weights[2529];
				12'd2530	: data <= weights[2530];
				12'd2531	: data <= weights[2531];
				12'd2532	: data <= weights[2532];
				12'd2533	: data <= weights[2533];
				12'd2534	: data <= weights[2534];
				12'd2535	: data <= weights[2535];
				12'd2536	: data <= weights[2536];
				12'd2537	: data <= weights[2537];
				12'd2538	: data <= weights[2538];
				12'd2539	: data <= weights[2539];
				12'd2540	: data <= weights[2540];
				12'd2541	: data <= weights[2541];
				12'd2542	: data <= weights[2542];
				12'd2543	: data <= weights[2543];
				12'd2544	: data <= weights[2544];
				12'd2545	: data <= weights[2545];
				12'd2546	: data <= weights[2546];
				12'd2547	: data <= weights[2547];
				12'd2548	: data <= weights[2548];
				12'd2549	: data <= weights[2549];
				12'd2550	: data <= weights[2550];
				12'd2551	: data <= weights[2551];
				12'd2552	: data <= weights[2552];
				12'd2553	: data <= weights[2553];
				12'd2554	: data <= weights[2554];
				12'd2555	: data <= weights[2555];
				12'd2556	: data <= weights[2556];
				12'd2557	: data <= weights[2557];
				12'd2558	: data <= weights[2558];
				12'd2559	: data <= weights[2559];
				12'd2560	: data <= weights[2560];
				12'd2561	: data <= weights[2561];
				12'd2562	: data <= weights[2562];
				12'd2563	: data <= weights[2563];
				12'd2564	: data <= weights[2564];
				12'd2565	: data <= weights[2565];
				12'd2566	: data <= weights[2566];
				12'd2567	: data <= weights[2567];
				12'd2568	: data <= weights[2568];
				12'd2569	: data <= weights[2569];
				12'd2570	: data <= weights[2570];
				12'd2571	: data <= weights[2571];
				12'd2572	: data <= weights[2572];
				12'd2573	: data <= weights[2573];
				12'd2574	: data <= weights[2574];
				12'd2575	: data <= weights[2575];
				12'd2576	: data <= weights[2576];
				12'd2577	: data <= weights[2577];
				12'd2578	: data <= weights[2578];
				12'd2579	: data <= weights[2579];
				12'd2580	: data <= weights[2580];
				12'd2581	: data <= weights[2581];
				12'd2582	: data <= weights[2582];
				12'd2583	: data <= weights[2583];
				12'd2584	: data <= weights[2584];
				12'd2585	: data <= weights[2585];
				12'd2586	: data <= weights[2586];
				12'd2587	: data <= weights[2587];
				12'd2588	: data <= weights[2588];
				12'd2589	: data <= weights[2589];
				12'd2590	: data <= weights[2590];
				12'd2591	: data <= weights[2591];
				12'd2592	: data <= weights[2592];
				12'd2593	: data <= weights[2593];
				12'd2594	: data <= weights[2594];
				12'd2595	: data <= weights[2595];
				12'd2596	: data <= weights[2596];
				12'd2597	: data <= weights[2597];
				12'd2598	: data <= weights[2598];
				12'd2599	: data <= weights[2599];
				12'd2600	: data <= weights[2600];
				12'd2601	: data <= weights[2601];
				12'd2602	: data <= weights[2602];
				12'd2603	: data <= weights[2603];
				12'd2604	: data <= weights[2604];
				12'd2605	: data <= weights[2605];
				12'd2606	: data <= weights[2606];
				12'd2607	: data <= weights[2607];
				12'd2608	: data <= weights[2608];
				12'd2609	: data <= weights[2609];
				12'd2610	: data <= weights[2610];
				12'd2611	: data <= weights[2611];
				12'd2612	: data <= weights[2612];
				12'd2613	: data <= weights[2613];
				12'd2614	: data <= weights[2614];
				12'd2615	: data <= weights[2615];
				12'd2616	: data <= weights[2616];
				12'd2617	: data <= weights[2617];
				12'd2618	: data <= weights[2618];
				12'd2619	: data <= weights[2619];
				12'd2620	: data <= weights[2620];
				12'd2621	: data <= weights[2621];
				12'd2622	: data <= weights[2622];
				12'd2623	: data <= weights[2623];
				12'd2624	: data <= weights[2624];
				12'd2625	: data <= weights[2625];
				12'd2626	: data <= weights[2626];
				12'd2627	: data <= weights[2627];
				12'd2628	: data <= weights[2628];
				12'd2629	: data <= weights[2629];
				12'd2630	: data <= weights[2630];
				12'd2631	: data <= weights[2631];
				12'd2632	: data <= weights[2632];
				12'd2633	: data <= weights[2633];
				12'd2634	: data <= weights[2634];
				12'd2635	: data <= weights[2635];
				12'd2636	: data <= weights[2636];
				12'd2637	: data <= weights[2637];
				12'd2638	: data <= weights[2638];
				12'd2639	: data <= weights[2639];
				12'd2640	: data <= weights[2640];
				12'd2641	: data <= weights[2641];
				12'd2642	: data <= weights[2642];
				12'd2643	: data <= weights[2643];
				12'd2644	: data <= weights[2644];
				12'd2645	: data <= weights[2645];
				12'd2646	: data <= weights[2646];
				12'd2647	: data <= weights[2647];
				12'd2648	: data <= weights[2648];
				12'd2649	: data <= weights[2649];
				12'd2650	: data <= weights[2650];
				12'd2651	: data <= weights[2651];
				12'd2652	: data <= weights[2652];
				12'd2653	: data <= weights[2653];
				12'd2654	: data <= weights[2654];
				12'd2655	: data <= weights[2655];
				12'd2656	: data <= weights[2656];
				12'd2657	: data <= weights[2657];
				12'd2658	: data <= weights[2658];
				12'd2659	: data <= weights[2659];
				12'd2660	: data <= weights[2660];
				12'd2661	: data <= weights[2661];
				12'd2662	: data <= weights[2662];
				12'd2663	: data <= weights[2663];
				12'd2664	: data <= weights[2664];
				12'd2665	: data <= weights[2665];
				12'd2666	: data <= weights[2666];
				12'd2667	: data <= weights[2667];
				12'd2668	: data <= weights[2668];
				12'd2669	: data <= weights[2669];
				12'd2670	: data <= weights[2670];
				12'd2671	: data <= weights[2671];
				12'd2672	: data <= weights[2672];
				12'd2673	: data <= weights[2673];
				12'd2674	: data <= weights[2674];
				12'd2675	: data <= weights[2675];
				12'd2676	: data <= weights[2676];
				12'd2677	: data <= weights[2677];
				12'd2678	: data <= weights[2678];
				12'd2679	: data <= weights[2679];
				12'd2680	: data <= weights[2680];
				12'd2681	: data <= weights[2681];
				12'd2682	: data <= weights[2682];
				12'd2683	: data <= weights[2683];
				12'd2684	: data <= weights[2684];
				12'd2685	: data <= weights[2685];
				12'd2686	: data <= weights[2686];
				12'd2687	: data <= weights[2687];
				12'd2688	: data <= weights[2688];
				12'd2689	: data <= weights[2689];
				12'd2690	: data <= weights[2690];
				12'd2691	: data <= weights[2691];
				12'd2692	: data <= weights[2692];
				12'd2693	: data <= weights[2693];
				12'd2694	: data <= weights[2694];
				12'd2695	: data <= weights[2695];
				12'd2696	: data <= weights[2696];
				12'd2697	: data <= weights[2697];
				12'd2698	: data <= weights[2698];
				12'd2699	: data <= weights[2699];
				12'd2700	: data <= weights[2700];
				12'd2701	: data <= weights[2701];
				12'd2702	: data <= weights[2702];
				12'd2703	: data <= weights[2703];
				12'd2704	: data <= weights[2704];
				12'd2705	: data <= weights[2705];
				12'd2706	: data <= weights[2706];
				12'd2707	: data <= weights[2707];
				12'd2708	: data <= weights[2708];
				12'd2709	: data <= weights[2709];
				12'd2710	: data <= weights[2710];
				12'd2711	: data <= weights[2711];
				12'd2712	: data <= weights[2712];
				12'd2713	: data <= weights[2713];
				12'd2714	: data <= weights[2714];
				12'd2715	: data <= weights[2715];
				12'd2716	: data <= weights[2716];
				12'd2717	: data <= weights[2717];
				12'd2718	: data <= weights[2718];
				12'd2719	: data <= weights[2719];
				12'd2720	: data <= weights[2720];
				12'd2721	: data <= weights[2721];
				12'd2722	: data <= weights[2722];
				12'd2723	: data <= weights[2723];
				12'd2724	: data <= weights[2724];
				12'd2725	: data <= weights[2725];
				12'd2726	: data <= weights[2726];
				12'd2727	: data <= weights[2727];
				12'd2728	: data <= weights[2728];
				12'd2729	: data <= weights[2729];
				12'd2730	: data <= weights[2730];
				12'd2731	: data <= weights[2731];
				12'd2732	: data <= weights[2732];
				12'd2733	: data <= weights[2733];
				12'd2734	: data <= weights[2734];
				12'd2735	: data <= weights[2735];
				12'd2736	: data <= weights[2736];
				12'd2737	: data <= weights[2737];
				12'd2738	: data <= weights[2738];
				12'd2739	: data <= weights[2739];
				12'd2740	: data <= weights[2740];
				12'd2741	: data <= weights[2741];
				12'd2742	: data <= weights[2742];
				12'd2743	: data <= weights[2743];
				12'd2744	: data <= weights[2744];
				12'd2745	: data <= weights[2745];
				12'd2746	: data <= weights[2746];
				12'd2747	: data <= weights[2747];
				12'd2748	: data <= weights[2748];
				12'd2749	: data <= weights[2749];
				12'd2750	: data <= weights[2750];
				12'd2751	: data <= weights[2751];
				12'd2752	: data <= weights[2752];
				12'd2753	: data <= weights[2753];
				12'd2754	: data <= weights[2754];
				12'd2755	: data <= weights[2755];
				12'd2756	: data <= weights[2756];
				12'd2757	: data <= weights[2757];
				12'd2758	: data <= weights[2758];
				12'd2759	: data <= weights[2759];
				12'd2760	: data <= weights[2760];
				12'd2761	: data <= weights[2761];
				12'd2762	: data <= weights[2762];
				12'd2763	: data <= weights[2763];
				12'd2764	: data <= weights[2764];
				12'd2765	: data <= weights[2765];
				12'd2766	: data <= weights[2766];
				12'd2767	: data <= weights[2767];
				12'd2768	: data <= weights[2768];
				12'd2769	: data <= weights[2769];
				12'd2770	: data <= weights[2770];
				12'd2771	: data <= weights[2771];
				12'd2772	: data <= weights[2772];
				12'd2773	: data <= weights[2773];
				12'd2774	: data <= weights[2774];
				12'd2775	: data <= weights[2775];
				12'd2776	: data <= weights[2776];
				12'd2777	: data <= weights[2777];
				12'd2778	: data <= weights[2778];
				12'd2779	: data <= weights[2779];
				12'd2780	: data <= weights[2780];
				12'd2781	: data <= weights[2781];
				12'd2782	: data <= weights[2782];
				12'd2783	: data <= weights[2783];
				12'd2784	: data <= weights[2784];
				12'd2785	: data <= weights[2785];
				12'd2786	: data <= weights[2786];
				12'd2787	: data <= weights[2787];
				12'd2788	: data <= weights[2788];
				12'd2789	: data <= weights[2789];
				12'd2790	: data <= weights[2790];
				12'd2791	: data <= weights[2791];
				12'd2792	: data <= weights[2792];
				12'd2793	: data <= weights[2793];
				12'd2794	: data <= weights[2794];
				12'd2795	: data <= weights[2795];
				12'd2796	: data <= weights[2796];
				12'd2797	: data <= weights[2797];
				12'd2798	: data <= weights[2798];
				12'd2799	: data <= weights[2799];
				12'd2800	: data <= weights[2800];
				12'd2801	: data <= weights[2801];
				12'd2802	: data <= weights[2802];
				12'd2803	: data <= weights[2803];
				12'd2804	: data <= weights[2804];
				12'd2805	: data <= weights[2805];
				12'd2806	: data <= weights[2806];
				12'd2807	: data <= weights[2807];
				12'd2808	: data <= weights[2808];
				12'd2809	: data <= weights[2809];
				12'd2810	: data <= weights[2810];
				12'd2811	: data <= weights[2811];
				12'd2812	: data <= weights[2812];
				12'd2813	: data <= weights[2813];
				12'd2814	: data <= weights[2814];
				12'd2815	: data <= weights[2815];
				12'd2816	: data <= weights[2816];
				12'd2817	: data <= weights[2817];
				12'd2818	: data <= weights[2818];
				12'd2819	: data <= weights[2819];
				12'd2820	: data <= weights[2820];
				12'd2821	: data <= weights[2821];
				12'd2822	: data <= weights[2822];
				12'd2823	: data <= weights[2823];
				12'd2824	: data <= weights[2824];
				12'd2825	: data <= weights[2825];
				12'd2826	: data <= weights[2826];
				12'd2827	: data <= weights[2827];
				12'd2828	: data <= weights[2828];
				12'd2829	: data <= weights[2829];
				12'd2830	: data <= weights[2830];
				12'd2831	: data <= weights[2831];
				12'd2832	: data <= weights[2832];
				12'd2833	: data <= weights[2833];
				12'd2834	: data <= weights[2834];
				12'd2835	: data <= weights[2835];
				12'd2836	: data <= weights[2836];
				12'd2837	: data <= weights[2837];
				12'd2838	: data <= weights[2838];
				12'd2839	: data <= weights[2839];
				12'd2840	: data <= weights[2840];
				12'd2841	: data <= weights[2841];
				12'd2842	: data <= weights[2842];
				12'd2843	: data <= weights[2843];
				12'd2844	: data <= weights[2844];
				12'd2845	: data <= weights[2845];
				12'd2846	: data <= weights[2846];
				12'd2847	: data <= weights[2847];
				12'd2848	: data <= weights[2848];
				12'd2849	: data <= weights[2849];
				12'd2850	: data <= weights[2850];
				12'd2851	: data <= weights[2851];
				12'd2852	: data <= weights[2852];
				12'd2853	: data <= weights[2853];
				12'd2854	: data <= weights[2854];
				12'd2855	: data <= weights[2855];
				12'd2856	: data <= weights[2856];
				12'd2857	: data <= weights[2857];
				12'd2858	: data <= weights[2858];
				12'd2859	: data <= weights[2859];
				12'd2860	: data <= weights[2860];
				12'd2861	: data <= weights[2861];
				12'd2862	: data <= weights[2862];
				12'd2863	: data <= weights[2863];
				12'd2864	: data <= weights[2864];
				12'd2865	: data <= weights[2865];
				12'd2866	: data <= weights[2866];
				12'd2867	: data <= weights[2867];
				12'd2868	: data <= weights[2868];
				12'd2869	: data <= weights[2869];
				12'd2870	: data <= weights[2870];
				12'd2871	: data <= weights[2871];
				12'd2872	: data <= weights[2872];
				12'd2873	: data <= weights[2873];
				12'd2874	: data <= weights[2874];
				12'd2875	: data <= weights[2875];
				12'd2876	: data <= weights[2876];
				12'd2877	: data <= weights[2877];
				12'd2878	: data <= weights[2878];
				12'd2879	: data <= weights[2879];
				12'd2880	: data <= weights[2880];
				12'd2881	: data <= weights[2881];
				12'd2882	: data <= weights[2882];
				12'd2883	: data <= weights[2883];
				12'd2884	: data <= weights[2884];
				12'd2885	: data <= weights[2885];
				12'd2886	: data <= weights[2886];
				12'd2887	: data <= weights[2887];
				12'd2888	: data <= weights[2888];
				12'd2889	: data <= weights[2889];
				12'd2890	: data <= weights[2890];
				12'd2891	: data <= weights[2891];
				12'd2892	: data <= weights[2892];
				12'd2893	: data <= weights[2893];
				12'd2894	: data <= weights[2894];
				12'd2895	: data <= weights[2895];
				12'd2896	: data <= weights[2896];
				12'd2897	: data <= weights[2897];
				12'd2898	: data <= weights[2898];
				12'd2899	: data <= weights[2899];
				12'd2900	: data <= weights[2900];
				12'd2901	: data <= weights[2901];
				12'd2902	: data <= weights[2902];
				12'd2903	: data <= weights[2903];
				12'd2904	: data <= weights[2904];
				12'd2905	: data <= weights[2905];
				12'd2906	: data <= weights[2906];
				12'd2907	: data <= weights[2907];
				12'd2908	: data <= weights[2908];
				12'd2909	: data <= weights[2909];
				12'd2910	: data <= weights[2910];
				12'd2911	: data <= weights[2911];
				12'd2912	: data <= weights[2912];
				12'd2913	: data <= weights[2913];
				12'd2914	: data <= weights[2914];
				12'd2915	: data <= weights[2915];
				12'd2916	: data <= weights[2916];
				12'd2917	: data <= weights[2917];
				12'd2918	: data <= weights[2918];
				12'd2919	: data <= weights[2919];
				12'd2920	: data <= weights[2920];
				12'd2921	: data <= weights[2921];
				12'd2922	: data <= weights[2922];
				12'd2923	: data <= weights[2923];
				12'd2924	: data <= weights[2924];
				12'd2925	: data <= weights[2925];
				12'd2926	: data <= weights[2926];
				12'd2927	: data <= weights[2927];
				12'd2928	: data <= weights[2928];
				12'd2929	: data <= weights[2929];
				12'd2930	: data <= weights[2930];
				12'd2931	: data <= weights[2931];
				12'd2932	: data <= weights[2932];
				12'd2933	: data <= weights[2933];
				12'd2934	: data <= weights[2934];
				12'd2935	: data <= weights[2935];
				12'd2936	: data <= weights[2936];
				12'd2937	: data <= weights[2937];
				12'd2938	: data <= weights[2938];
				12'd2939	: data <= weights[2939];
				12'd2940	: data <= weights[2940];
				12'd2941	: data <= weights[2941];
				12'd2942	: data <= weights[2942];
				12'd2943	: data <= weights[2943];
				12'd2944	: data <= weights[2944];
				12'd2945	: data <= weights[2945];
				12'd2946	: data <= weights[2946];
				12'd2947	: data <= weights[2947];
				12'd2948	: data <= weights[2948];
				12'd2949	: data <= weights[2949];
				12'd2950	: data <= weights[2950];
				12'd2951	: data <= weights[2951];
				12'd2952	: data <= weights[2952];
				12'd2953	: data <= weights[2953];
				12'd2954	: data <= weights[2954];
				12'd2955	: data <= weights[2955];
				12'd2956	: data <= weights[2956];
				12'd2957	: data <= weights[2957];
				12'd2958	: data <= weights[2958];
				12'd2959	: data <= weights[2959];
				12'd2960	: data <= weights[2960];
				12'd2961	: data <= weights[2961];
				12'd2962	: data <= weights[2962];
				12'd2963	: data <= weights[2963];
				12'd2964	: data <= weights[2964];
				12'd2965	: data <= weights[2965];
				12'd2966	: data <= weights[2966];
				12'd2967	: data <= weights[2967];
				12'd2968	: data <= weights[2968];
				12'd2969	: data <= weights[2969];
				12'd2970	: data <= weights[2970];
				12'd2971	: data <= weights[2971];
				12'd2972	: data <= weights[2972];
				12'd2973	: data <= weights[2973];
				12'd2974	: data <= weights[2974];
				12'd2975	: data <= weights[2975];
				12'd2976	: data <= weights[2976];
				12'd2977	: data <= weights[2977];
				12'd2978	: data <= weights[2978];
				12'd2979	: data <= weights[2979];
				12'd2980	: data <= weights[2980];
				12'd2981	: data <= weights[2981];
				12'd2982	: data <= weights[2982];
				12'd2983	: data <= weights[2983];
				12'd2984	: data <= weights[2984];
				12'd2985	: data <= weights[2985];
				12'd2986	: data <= weights[2986];
				12'd2987	: data <= weights[2987];
				12'd2988	: data <= weights[2988];
				12'd2989	: data <= weights[2989];
				12'd2990	: data <= weights[2990];
				12'd2991	: data <= weights[2991];
				12'd2992	: data <= weights[2992];
				12'd2993	: data <= weights[2993];
				12'd2994	: data <= weights[2994];
				12'd2995	: data <= weights[2995];
				12'd2996	: data <= weights[2996];
				12'd2997	: data <= weights[2997];
				12'd2998	: data <= weights[2998];
				12'd2999	: data <= weights[2999];
				12'd3000	: data <= weights[3000];
				12'd3001	: data <= weights[3001];
				12'd3002	: data <= weights[3002];
				12'd3003	: data <= weights[3003];
				12'd3004	: data <= weights[3004];
				12'd3005	: data <= weights[3005];
				12'd3006	: data <= weights[3006];
				12'd3007	: data <= weights[3007];
				12'd3008	: data <= weights[3008];
				12'd3009	: data <= weights[3009];
				12'd3010	: data <= weights[3010];
				12'd3011	: data <= weights[3011];
				12'd3012	: data <= weights[3012];
				12'd3013	: data <= weights[3013];
				12'd3014	: data <= weights[3014];
				12'd3015	: data <= weights[3015];
				12'd3016	: data <= weights[3016];
				12'd3017	: data <= weights[3017];
				12'd3018	: data <= weights[3018];
				12'd3019	: data <= weights[3019];
				12'd3020	: data <= weights[3020];
				12'd3021	: data <= weights[3021];
				12'd3022	: data <= weights[3022];
				12'd3023	: data <= weights[3023];
				12'd3024	: data <= weights[3024];
				12'd3025	: data <= weights[3025];
				12'd3026	: data <= weights[3026];
				12'd3027	: data <= weights[3027];
				12'd3028	: data <= weights[3028];
				12'd3029	: data <= weights[3029];
				12'd3030	: data <= weights[3030];
				12'd3031	: data <= weights[3031];
				12'd3032	: data <= weights[3032];
				12'd3033	: data <= weights[3033];
				12'd3034	: data <= weights[3034];
				12'd3035	: data <= weights[3035];
				12'd3036	: data <= weights[3036];
				12'd3037	: data <= weights[3037];
				12'd3038	: data <= weights[3038];
				12'd3039	: data <= weights[3039];
				12'd3040	: data <= weights[3040];
				12'd3041	: data <= weights[3041];
				12'd3042	: data <= weights[3042];
				12'd3043	: data <= weights[3043];
				12'd3044	: data <= weights[3044];
				12'd3045	: data <= weights[3045];
				12'd3046	: data <= weights[3046];
				12'd3047	: data <= weights[3047];
				12'd3048	: data <= weights[3048];
				12'd3049	: data <= weights[3049];
				12'd3050	: data <= weights[3050];
				12'd3051	: data <= weights[3051];
				12'd3052	: data <= weights[3052];
				12'd3053	: data <= weights[3053];
				12'd3054	: data <= weights[3054];
				12'd3055	: data <= weights[3055];
				12'd3056	: data <= weights[3056];
				12'd3057	: data <= weights[3057];
				12'd3058	: data <= weights[3058];
				12'd3059	: data <= weights[3059];
				12'd3060	: data <= weights[3060];
				12'd3061	: data <= weights[3061];
				12'd3062	: data <= weights[3062];
				12'd3063	: data <= weights[3063];
				12'd3064	: data <= weights[3064];
				12'd3065	: data <= weights[3065];
				12'd3066	: data <= weights[3066];
				12'd3067	: data <= weights[3067];
				12'd3068	: data <= weights[3068];
				12'd3069	: data <= weights[3069];
				12'd3070	: data <= weights[3070];
				12'd3071	: data <= weights[3071];
				12'd3072	: data <= weights[3072];
				12'd3073	: data <= weights[3073];
				12'd3074	: data <= weights[3074];
				12'd3075	: data <= weights[3075];
				12'd3076	: data <= weights[3076];
				12'd3077	: data <= weights[3077];
				12'd3078	: data <= weights[3078];
				12'd3079	: data <= weights[3079];
				12'd3080	: data <= weights[3080];
				12'd3081	: data <= weights[3081];
				12'd3082	: data <= weights[3082];
				12'd3083	: data <= weights[3083];
				12'd3084	: data <= weights[3084];
				12'd3085	: data <= weights[3085];
				12'd3086	: data <= weights[3086];
				12'd3087	: data <= weights[3087];
				12'd3088	: data <= weights[3088];
				12'd3089	: data <= weights[3089];
				12'd3090	: data <= weights[3090];
				12'd3091	: data <= weights[3091];
				12'd3092	: data <= weights[3092];
				12'd3093	: data <= weights[3093];
				12'd3094	: data <= weights[3094];
				12'd3095	: data <= weights[3095];
				12'd3096	: data <= weights[3096];
				12'd3097	: data <= weights[3097];
				12'd3098	: data <= weights[3098];
				12'd3099	: data <= weights[3099];
				12'd3100	: data <= weights[3100];
				12'd3101	: data <= weights[3101];
				12'd3102	: data <= weights[3102];
				12'd3103	: data <= weights[3103];
				12'd3104	: data <= weights[3104];
				12'd3105	: data <= weights[3105];
				12'd3106	: data <= weights[3106];
				12'd3107	: data <= weights[3107];
				12'd3108	: data <= weights[3108];
				12'd3109	: data <= weights[3109];
				12'd3110	: data <= weights[3110];
				12'd3111	: data <= weights[3111];
				12'd3112	: data <= weights[3112];
				12'd3113	: data <= weights[3113];
				12'd3114	: data <= weights[3114];
				12'd3115	: data <= weights[3115];
				12'd3116	: data <= weights[3116];
				12'd3117	: data <= weights[3117];
				12'd3118	: data <= weights[3118];
				12'd3119	: data <= weights[3119];
				12'd3120	: data <= weights[3120];
				12'd3121	: data <= weights[3121];
				12'd3122	: data <= weights[3122];
				12'd3123	: data <= weights[3123];
				12'd3124	: data <= weights[3124];
				12'd3125	: data <= weights[3125];
				12'd3126	: data <= weights[3126];
				12'd3127	: data <= weights[3127];
				12'd3128	: data <= weights[3128];
				12'd3129	: data <= weights[3129];
				12'd3130	: data <= weights[3130];
				12'd3131	: data <= weights[3131];
				12'd3132	: data <= weights[3132];
				12'd3133	: data <= weights[3133];
				12'd3134	: data <= weights[3134];
				12'd3135	: data <= weights[3135];
				12'd3136	: data <= weights[3136];
				12'd3137	: data <= weights[3137];
				12'd3138	: data <= weights[3138];
				12'd3139	: data <= weights[3139];
				12'd3140	: data <= weights[3140];
				12'd3141	: data <= weights[3141];
				12'd3142	: data <= weights[3142];
				12'd3143	: data <= weights[3143];
				12'd3144	: data <= weights[3144];
				12'd3145	: data <= weights[3145];
				12'd3146	: data <= weights[3146];
				12'd3147	: data <= weights[3147];
				12'd3148	: data <= weights[3148];
				12'd3149	: data <= weights[3149];
				12'd3150	: data <= weights[3150];
				12'd3151	: data <= weights[3151];
				12'd3152	: data <= weights[3152];
				12'd3153	: data <= weights[3153];
				12'd3154	: data <= weights[3154];
				12'd3155	: data <= weights[3155];
				12'd3156	: data <= weights[3156];
				12'd3157	: data <= weights[3157];
				12'd3158	: data <= weights[3158];
				12'd3159	: data <= weights[3159];
				12'd3160	: data <= weights[3160];
				12'd3161	: data <= weights[3161];
				12'd3162	: data <= weights[3162];
				12'd3163	: data <= weights[3163];
				12'd3164	: data <= weights[3164];
				12'd3165	: data <= weights[3165];
				12'd3166	: data <= weights[3166];
				12'd3167	: data <= weights[3167];
				12'd3168	: data <= weights[3168];
				12'd3169	: data <= weights[3169];
				12'd3170	: data <= weights[3170];
				12'd3171	: data <= weights[3171];
				12'd3172	: data <= weights[3172];
				12'd3173	: data <= weights[3173];
				12'd3174	: data <= weights[3174];
				12'd3175	: data <= weights[3175];
				12'd3176	: data <= weights[3176];
				12'd3177	: data <= weights[3177];
				12'd3178	: data <= weights[3178];
				12'd3179	: data <= weights[3179];
				12'd3180	: data <= weights[3180];
				12'd3181	: data <= weights[3181];
				12'd3182	: data <= weights[3182];
				12'd3183	: data <= weights[3183];
				12'd3184	: data <= weights[3184];
				12'd3185	: data <= weights[3185];
				12'd3186	: data <= weights[3186];
				12'd3187	: data <= weights[3187];
				12'd3188	: data <= weights[3188];
				12'd3189	: data <= weights[3189];
				12'd3190	: data <= weights[3190];
				12'd3191	: data <= weights[3191];
				12'd3192	: data <= weights[3192];
				12'd3193	: data <= weights[3193];
				12'd3194	: data <= weights[3194];
				12'd3195	: data <= weights[3195];
				12'd3196	: data <= weights[3196];
				12'd3197	: data <= weights[3197];
				12'd3198	: data <= weights[3198];
				12'd3199	: data <= weights[3199];
				12'd3200	: data <= weights[3200];
				12'd3201	: data <= weights[3201];
				12'd3202	: data <= weights[3202];
				12'd3203	: data <= weights[3203];
				12'd3204	: data <= weights[3204];
				12'd3205	: data <= weights[3205];
				12'd3206	: data <= weights[3206];
				12'd3207	: data <= weights[3207];
				12'd3208	: data <= weights[3208];
				12'd3209	: data <= weights[3209];
				12'd3210	: data <= weights[3210];
				12'd3211	: data <= weights[3211];
				12'd3212	: data <= weights[3212];
				12'd3213	: data <= weights[3213];
				12'd3214	: data <= weights[3214];
				12'd3215	: data <= weights[3215];
				12'd3216	: data <= weights[3216];
				12'd3217	: data <= weights[3217];
				12'd3218	: data <= weights[3218];
				12'd3219	: data <= weights[3219];
				12'd3220	: data <= weights[3220];
				12'd3221	: data <= weights[3221];
				12'd3222	: data <= weights[3222];
				12'd3223	: data <= weights[3223];
				12'd3224	: data <= weights[3224];
				12'd3225	: data <= weights[3225];
				12'd3226	: data <= weights[3226];
				12'd3227	: data <= weights[3227];
				12'd3228	: data <= weights[3228];
				12'd3229	: data <= weights[3229];
				12'd3230	: data <= weights[3230];
				12'd3231	: data <= weights[3231];
				12'd3232	: data <= weights[3232];
				12'd3233	: data <= weights[3233];
				12'd3234	: data <= weights[3234];
				12'd3235	: data <= weights[3235];
				12'd3236	: data <= weights[3236];
				12'd3237	: data <= weights[3237];
				12'd3238	: data <= weights[3238];
				12'd3239	: data <= weights[3239];
				12'd3240	: data <= weights[3240];
				12'd3241	: data <= weights[3241];
				12'd3242	: data <= weights[3242];
				12'd3243	: data <= weights[3243];
				12'd3244	: data <= weights[3244];
				12'd3245	: data <= weights[3245];
				12'd3246	: data <= weights[3246];
				12'd3247	: data <= weights[3247];
				12'd3248	: data <= weights[3248];
				12'd3249	: data <= weights[3249];
				12'd3250	: data <= weights[3250];
				12'd3251	: data <= weights[3251];
				12'd3252	: data <= weights[3252];
				12'd3253	: data <= weights[3253];
				12'd3254	: data <= weights[3254];
				12'd3255	: data <= weights[3255];
				12'd3256	: data <= weights[3256];
				12'd3257	: data <= weights[3257];
				12'd3258	: data <= weights[3258];
				12'd3259	: data <= weights[3259];
				12'd3260	: data <= weights[3260];
				12'd3261	: data <= weights[3261];
				12'd3262	: data <= weights[3262];
				12'd3263	: data <= weights[3263];
				12'd3264	: data <= weights[3264];
				12'd3265	: data <= weights[3265];
				12'd3266	: data <= weights[3266];
				12'd3267	: data <= weights[3267];
				12'd3268	: data <= weights[3268];
				12'd3269	: data <= weights[3269];
				12'd3270	: data <= weights[3270];
				12'd3271	: data <= weights[3271];
				12'd3272	: data <= weights[3272];
				12'd3273	: data <= weights[3273];
				12'd3274	: data <= weights[3274];
				12'd3275	: data <= weights[3275];
				12'd3276	: data <= weights[3276];
				12'd3277	: data <= weights[3277];
				12'd3278	: data <= weights[3278];
				12'd3279	: data <= weights[3279];
				12'd3280	: data <= weights[3280];
				12'd3281	: data <= weights[3281];
				12'd3282	: data <= weights[3282];
				12'd3283	: data <= weights[3283];
				12'd3284	: data <= weights[3284];
				12'd3285	: data <= weights[3285];
				12'd3286	: data <= weights[3286];
				12'd3287	: data <= weights[3287];
				12'd3288	: data <= weights[3288];
				12'd3289	: data <= weights[3289];
				12'd3290	: data <= weights[3290];
				12'd3291	: data <= weights[3291];
				12'd3292	: data <= weights[3292];
				12'd3293	: data <= weights[3293];
				12'd3294	: data <= weights[3294];
				12'd3295	: data <= weights[3295];
				12'd3296	: data <= weights[3296];
				12'd3297	: data <= weights[3297];
				12'd3298	: data <= weights[3298];
				12'd3299	: data <= weights[3299];
				12'd3300	: data <= weights[3300];
				12'd3301	: data <= weights[3301];
				12'd3302	: data <= weights[3302];
				12'd3303	: data <= weights[3303];
				12'd3304	: data <= weights[3304];
				12'd3305	: data <= weights[3305];
				12'd3306	: data <= weights[3306];
				12'd3307	: data <= weights[3307];
				12'd3308	: data <= weights[3308];
				12'd3309	: data <= weights[3309];
				12'd3310	: data <= weights[3310];
				12'd3311	: data <= weights[3311];
				12'd3312	: data <= weights[3312];
				12'd3313	: data <= weights[3313];
				12'd3314	: data <= weights[3314];
				12'd3315	: data <= weights[3315];
				12'd3316	: data <= weights[3316];
				12'd3317	: data <= weights[3317];
				12'd3318	: data <= weights[3318];
				12'd3319	: data <= weights[3319];
				12'd3320	: data <= weights[3320];
				12'd3321	: data <= weights[3321];
				12'd3322	: data <= weights[3322];
				12'd3323	: data <= weights[3323];
				12'd3324	: data <= weights[3324];
				12'd3325	: data <= weights[3325];
				12'd3326	: data <= weights[3326];
				12'd3327	: data <= weights[3327];
				12'd3328	: data <= weights[3328];
				12'd3329	: data <= weights[3329];
				12'd3330	: data <= weights[3330];
				12'd3331	: data <= weights[3331];
				12'd3332	: data <= weights[3332];
				12'd3333	: data <= weights[3333];
				12'd3334	: data <= weights[3334];
				12'd3335	: data <= weights[3335];
				12'd3336	: data <= weights[3336];
				12'd3337	: data <= weights[3337];
				12'd3338	: data <= weights[3338];
				12'd3339	: data <= weights[3339];
				12'd3340	: data <= weights[3340];
				12'd3341	: data <= weights[3341];
				12'd3342	: data <= weights[3342];
				12'd3343	: data <= weights[3343];
				12'd3344	: data <= weights[3344];
				12'd3345	: data <= weights[3345];
				12'd3346	: data <= weights[3346];
				12'd3347	: data <= weights[3347];
				12'd3348	: data <= weights[3348];
				12'd3349	: data <= weights[3349];
				12'd3350	: data <= weights[3350];
				12'd3351	: data <= weights[3351];
				12'd3352	: data <= weights[3352];
				12'd3353	: data <= weights[3353];
				12'd3354	: data <= weights[3354];
				12'd3355	: data <= weights[3355];
				12'd3356	: data <= weights[3356];
				12'd3357	: data <= weights[3357];
				12'd3358	: data <= weights[3358];
				12'd3359	: data <= weights[3359];
				12'd3360	: data <= weights[3360];
				12'd3361	: data <= weights[3361];
				12'd3362	: data <= weights[3362];
				12'd3363	: data <= weights[3363];
				12'd3364	: data <= weights[3364];
				12'd3365	: data <= weights[3365];
				12'd3366	: data <= weights[3366];
				12'd3367	: data <= weights[3367];
				12'd3368	: data <= weights[3368];
				12'd3369	: data <= weights[3369];
				12'd3370	: data <= weights[3370];
				12'd3371	: data <= weights[3371];
				12'd3372	: data <= weights[3372];
				12'd3373	: data <= weights[3373];
				12'd3374	: data <= weights[3374];
				12'd3375	: data <= weights[3375];
				12'd3376	: data <= weights[3376];
				12'd3377	: data <= weights[3377];
				12'd3378	: data <= weights[3378];
				12'd3379	: data <= weights[3379];
				12'd3380	: data <= weights[3380];
				12'd3381	: data <= weights[3381];
				12'd3382	: data <= weights[3382];
				12'd3383	: data <= weights[3383];
				12'd3384	: data <= weights[3384];
				12'd3385	: data <= weights[3385];
				12'd3386	: data <= weights[3386];
				12'd3387	: data <= weights[3387];
				12'd3388	: data <= weights[3388];
				12'd3389	: data <= weights[3389];
				12'd3390	: data <= weights[3390];
				12'd3391	: data <= weights[3391];
				12'd3392	: data <= weights[3392];
				12'd3393	: data <= weights[3393];
				12'd3394	: data <= weights[3394];
				12'd3395	: data <= weights[3395];
				12'd3396	: data <= weights[3396];
				12'd3397	: data <= weights[3397];
				12'd3398	: data <= weights[3398];
				12'd3399	: data <= weights[3399];
				12'd3400	: data <= weights[3400];
				12'd3401	: data <= weights[3401];
				12'd3402	: data <= weights[3402];
				12'd3403	: data <= weights[3403];
				12'd3404	: data <= weights[3404];
				12'd3405	: data <= weights[3405];
				12'd3406	: data <= weights[3406];
				12'd3407	: data <= weights[3407];
				12'd3408	: data <= weights[3408];
				12'd3409	: data <= weights[3409];
				12'd3410	: data <= weights[3410];
				12'd3411	: data <= weights[3411];
				12'd3412	: data <= weights[3412];
				12'd3413	: data <= weights[3413];
				12'd3414	: data <= weights[3414];
				12'd3415	: data <= weights[3415];
				12'd3416	: data <= weights[3416];
				12'd3417	: data <= weights[3417];
				12'd3418	: data <= weights[3418];
				12'd3419	: data <= weights[3419];
				12'd3420	: data <= weights[3420];
				12'd3421	: data <= weights[3421];
				12'd3422	: data <= weights[3422];
				12'd3423	: data <= weights[3423];
				12'd3424	: data <= weights[3424];
				12'd3425	: data <= weights[3425];
				12'd3426	: data <= weights[3426];
				12'd3427	: data <= weights[3427];
				12'd3428	: data <= weights[3428];
				12'd3429	: data <= weights[3429];
				12'd3430	: data <= weights[3430];
				12'd3431	: data <= weights[3431];
				12'd3432	: data <= weights[3432];
				12'd3433	: data <= weights[3433];
				12'd3434	: data <= weights[3434];
				12'd3435	: data <= weights[3435];
				12'd3436	: data <= weights[3436];
				12'd3437	: data <= weights[3437];
				12'd3438	: data <= weights[3438];
				12'd3439	: data <= weights[3439];
				12'd3440	: data <= weights[3440];
				12'd3441	: data <= weights[3441];
				12'd3442	: data <= weights[3442];
				12'd3443	: data <= weights[3443];
				12'd3444	: data <= weights[3444];
				12'd3445	: data <= weights[3445];
				12'd3446	: data <= weights[3446];
				12'd3447	: data <= weights[3447];
				12'd3448	: data <= weights[3448];
				12'd3449	: data <= weights[3449];
				12'd3450	: data <= weights[3450];
				12'd3451	: data <= weights[3451];
				12'd3452	: data <= weights[3452];
				12'd3453	: data <= weights[3453];
				12'd3454	: data <= weights[3454];
				12'd3455	: data <= weights[3455];
				12'd3456	: data <= weights[3456];
				12'd3457	: data <= weights[3457];
				12'd3458	: data <= weights[3458];
				12'd3459	: data <= weights[3459];
				12'd3460	: data <= weights[3460];
				12'd3461	: data <= weights[3461];
				12'd3462	: data <= weights[3462];
				12'd3463	: data <= weights[3463];
				12'd3464	: data <= weights[3464];
				12'd3465	: data <= weights[3465];
				12'd3466	: data <= weights[3466];
				12'd3467	: data <= weights[3467];
				12'd3468	: data <= weights[3468];
				12'd3469	: data <= weights[3469];
				12'd3470	: data <= weights[3470];
				12'd3471	: data <= weights[3471];
				12'd3472	: data <= weights[3472];
				12'd3473	: data <= weights[3473];
				12'd3474	: data <= weights[3474];
				12'd3475	: data <= weights[3475];
				12'd3476	: data <= weights[3476];
				12'd3477	: data <= weights[3477];
				12'd3478	: data <= weights[3478];
				12'd3479	: data <= weights[3479];
				12'd3480	: data <= weights[3480];
				12'd3481	: data <= weights[3481];
				12'd3482	: data <= weights[3482];
				12'd3483	: data <= weights[3483];
				12'd3484	: data <= weights[3484];
				12'd3485	: data <= weights[3485];
				12'd3486	: data <= weights[3486];
				12'd3487	: data <= weights[3487];
				12'd3488	: data <= weights[3488];
				12'd3489	: data <= weights[3489];
				12'd3490	: data <= weights[3490];
				12'd3491	: data <= weights[3491];
				12'd3492	: data <= weights[3492];
				12'd3493	: data <= weights[3493];
				12'd3494	: data <= weights[3494];
				12'd3495	: data <= weights[3495];
				12'd3496	: data <= weights[3496];
				12'd3497	: data <= weights[3497];
				12'd3498	: data <= weights[3498];
				12'd3499	: data <= weights[3499];
				12'd3500	: data <= weights[3500];
				12'd3501	: data <= weights[3501];
				12'd3502	: data <= weights[3502];
				12'd3503	: data <= weights[3503];
				12'd3504	: data <= weights[3504];
				12'd3505	: data <= weights[3505];
				12'd3506	: data <= weights[3506];
				12'd3507	: data <= weights[3507];
				12'd3508	: data <= weights[3508];
				12'd3509	: data <= weights[3509];
				12'd3510	: data <= weights[3510];
				12'd3511	: data <= weights[3511];
				12'd3512	: data <= weights[3512];
				12'd3513	: data <= weights[3513];
				12'd3514	: data <= weights[3514];
				12'd3515	: data <= weights[3515];
				12'd3516	: data <= weights[3516];
				12'd3517	: data <= weights[3517];
				12'd3518	: data <= weights[3518];
				12'd3519	: data <= weights[3519];
				12'd3520	: data <= weights[3520];
				12'd3521	: data <= weights[3521];
				12'd3522	: data <= weights[3522];
				12'd3523	: data <= weights[3523];
				12'd3524	: data <= weights[3524];
				12'd3525	: data <= weights[3525];
				12'd3526	: data <= weights[3526];
				12'd3527	: data <= weights[3527];
				12'd3528	: data <= weights[3528];
				12'd3529	: data <= weights[3529];
				12'd3530	: data <= weights[3530];
				12'd3531	: data <= weights[3531];
				12'd3532	: data <= weights[3532];
				12'd3533	: data <= weights[3533];
				12'd3534	: data <= weights[3534];
				12'd3535	: data <= weights[3535];
				12'd3536	: data <= weights[3536];
				12'd3537	: data <= weights[3537];
				12'd3538	: data <= weights[3538];
				12'd3539	: data <= weights[3539];
				12'd3540	: data <= weights[3540];
				12'd3541	: data <= weights[3541];
				12'd3542	: data <= weights[3542];
				12'd3543	: data <= weights[3543];
				12'd3544	: data <= weights[3544];
				12'd3545	: data <= weights[3545];
				12'd3546	: data <= weights[3546];
				12'd3547	: data <= weights[3547];
				12'd3548	: data <= weights[3548];
				12'd3549	: data <= weights[3549];
				12'd3550	: data <= weights[3550];
				12'd3551	: data <= weights[3551];
				12'd3552	: data <= weights[3552];
				12'd3553	: data <= weights[3553];
				12'd3554	: data <= weights[3554];
				12'd3555	: data <= weights[3555];
				12'd3556	: data <= weights[3556];
				12'd3557	: data <= weights[3557];
				12'd3558	: data <= weights[3558];
				12'd3559	: data <= weights[3559];
				12'd3560	: data <= weights[3560];
				12'd3561	: data <= weights[3561];
				12'd3562	: data <= weights[3562];
				12'd3563	: data <= weights[3563];
				12'd3564	: data <= weights[3564];
				12'd3565	: data <= weights[3565];
				12'd3566	: data <= weights[3566];
				12'd3567	: data <= weights[3567];
				12'd3568	: data <= weights[3568];
				12'd3569	: data <= weights[3569];
				12'd3570	: data <= weights[3570];
				12'd3571	: data <= weights[3571];
				12'd3572	: data <= weights[3572];
				12'd3573	: data <= weights[3573];
				12'd3574	: data <= weights[3574];
				12'd3575	: data <= weights[3575];
				12'd3576	: data <= weights[3576];
				12'd3577	: data <= weights[3577];
				12'd3578	: data <= weights[3578];
				12'd3579	: data <= weights[3579];
				12'd3580	: data <= weights[3580];
				12'd3581	: data <= weights[3581];
				12'd3582	: data <= weights[3582];
				12'd3583	: data <= weights[3583];
				12'd3584	: data <= weights[3584];
				12'd3585	: data <= weights[3585];
				12'd3586	: data <= weights[3586];
				12'd3587	: data <= weights[3587];
				12'd3588	: data <= weights[3588];
				12'd3589	: data <= weights[3589];
				12'd3590	: data <= weights[3590];
				12'd3591	: data <= weights[3591];
				12'd3592	: data <= weights[3592];
				12'd3593	: data <= weights[3593];
				12'd3594	: data <= weights[3594];
				12'd3595	: data <= weights[3595];
				12'd3596	: data <= weights[3596];
				12'd3597	: data <= weights[3597];
				12'd3598	: data <= weights[3598];
				12'd3599	: data <= weights[3599];
				12'd3600	: data <= weights[3600];
				12'd3601	: data <= weights[3601];
				12'd3602	: data <= weights[3602];
				12'd3603	: data <= weights[3603];
				12'd3604	: data <= weights[3604];
				12'd3605	: data <= weights[3605];
				12'd3606	: data <= weights[3606];
				12'd3607	: data <= weights[3607];
				12'd3608	: data <= weights[3608];
				12'd3609	: data <= weights[3609];
				12'd3610	: data <= weights[3610];
				12'd3611	: data <= weights[3611];
				12'd3612	: data <= weights[3612];
				12'd3613	: data <= weights[3613];
				12'd3614	: data <= weights[3614];
				12'd3615	: data <= weights[3615];
				12'd3616	: data <= weights[3616];
				12'd3617	: data <= weights[3617];
				12'd3618	: data <= weights[3618];
				12'd3619	: data <= weights[3619];
				12'd3620	: data <= weights[3620];
				12'd3621	: data <= weights[3621];
				12'd3622	: data <= weights[3622];
				12'd3623	: data <= weights[3623];
				12'd3624	: data <= weights[3624];
				12'd3625	: data <= weights[3625];
				12'd3626	: data <= weights[3626];
				12'd3627	: data <= weights[3627];
				12'd3628	: data <= weights[3628];
				12'd3629	: data <= weights[3629];
				12'd3630	: data <= weights[3630];
				12'd3631	: data <= weights[3631];
				12'd3632	: data <= weights[3632];
				12'd3633	: data <= weights[3633];
				12'd3634	: data <= weights[3634];
				12'd3635	: data <= weights[3635];
				12'd3636	: data <= weights[3636];
				12'd3637	: data <= weights[3637];
				12'd3638	: data <= weights[3638];
				12'd3639	: data <= weights[3639];
				12'd3640	: data <= weights[3640];
				12'd3641	: data <= weights[3641];
				12'd3642	: data <= weights[3642];
				12'd3643	: data <= weights[3643];
				12'd3644	: data <= weights[3644];
				12'd3645	: data <= weights[3645];
				12'd3646	: data <= weights[3646];
				12'd3647	: data <= weights[3647];
				12'd3648	: data <= weights[3648];
				12'd3649	: data <= weights[3649];
				12'd3650	: data <= weights[3650];
				12'd3651	: data <= weights[3651];
				12'd3652	: data <= weights[3652];
				12'd3653	: data <= weights[3653];
				12'd3654	: data <= weights[3654];
				12'd3655	: data <= weights[3655];
				12'd3656	: data <= weights[3656];
				12'd3657	: data <= weights[3657];
				12'd3658	: data <= weights[3658];
				12'd3659	: data <= weights[3659];
				12'd3660	: data <= weights[3660];
				12'd3661	: data <= weights[3661];
				12'd3662	: data <= weights[3662];
				12'd3663	: data <= weights[3663];
				12'd3664	: data <= weights[3664];
				12'd3665	: data <= weights[3665];
				12'd3666	: data <= weights[3666];
				12'd3667	: data <= weights[3667];
				12'd3668	: data <= weights[3668];
				12'd3669	: data <= weights[3669];
				12'd3670	: data <= weights[3670];
				12'd3671	: data <= weights[3671];
				12'd3672	: data <= weights[3672];
				12'd3673	: data <= weights[3673];
				12'd3674	: data <= weights[3674];
				12'd3675	: data <= weights[3675];
				12'd3676	: data <= weights[3676];
				12'd3677	: data <= weights[3677];
				12'd3678	: data <= weights[3678];
				12'd3679	: data <= weights[3679];
				12'd3680	: data <= weights[3680];
				12'd3681	: data <= weights[3681];
				12'd3682	: data <= weights[3682];
				12'd3683	: data <= weights[3683];
				12'd3684	: data <= weights[3684];
				12'd3685	: data <= weights[3685];
				12'd3686	: data <= weights[3686];
				12'd3687	: data <= weights[3687];
				12'd3688	: data <= weights[3688];
				12'd3689	: data <= weights[3689];
				12'd3690	: data <= weights[3690];
				12'd3691	: data <= weights[3691];
				12'd3692	: data <= weights[3692];
				12'd3693	: data <= weights[3693];
				12'd3694	: data <= weights[3694];
				12'd3695	: data <= weights[3695];
				12'd3696	: data <= weights[3696];
				12'd3697	: data <= weights[3697];
				12'd3698	: data <= weights[3698];
				12'd3699	: data <= weights[3699];
				12'd3700	: data <= weights[3700];
				12'd3701	: data <= weights[3701];
				12'd3702	: data <= weights[3702];
				12'd3703	: data <= weights[3703];
				12'd3704	: data <= weights[3704];
				12'd3705	: data <= weights[3705];
				12'd3706	: data <= weights[3706];
				12'd3707	: data <= weights[3707];
				12'd3708	: data <= weights[3708];
				12'd3709	: data <= weights[3709];
				12'd3710	: data <= weights[3710];
				12'd3711	: data <= weights[3711];
				12'd3712	: data <= weights[3712];
				12'd3713	: data <= weights[3713];
				12'd3714	: data <= weights[3714];
				12'd3715	: data <= weights[3715];
				12'd3716	: data <= weights[3716];
				12'd3717	: data <= weights[3717];
				12'd3718	: data <= weights[3718];
				12'd3719	: data <= weights[3719];
				12'd3720	: data <= weights[3720];
				12'd3721	: data <= weights[3721];
				12'd3722	: data <= weights[3722];
				12'd3723	: data <= weights[3723];
				12'd3724	: data <= weights[3724];
				12'd3725	: data <= weights[3725];
				12'd3726	: data <= weights[3726];
				12'd3727	: data <= weights[3727];
				12'd3728	: data <= weights[3728];
				12'd3729	: data <= weights[3729];
				12'd3730	: data <= weights[3730];
				12'd3731	: data <= weights[3731];
				12'd3732	: data <= weights[3732];
				12'd3733	: data <= weights[3733];
				12'd3734	: data <= weights[3734];
				12'd3735	: data <= weights[3735];
				12'd3736	: data <= weights[3736];
				12'd3737	: data <= weights[3737];
				12'd3738	: data <= weights[3738];
				12'd3739	: data <= weights[3739];
				12'd3740	: data <= weights[3740];
				12'd3741	: data <= weights[3741];
				12'd3742	: data <= weights[3742];
				12'd3743	: data <= weights[3743];
				12'd3744	: data <= weights[3744];
				12'd3745	: data <= weights[3745];
				12'd3746	: data <= weights[3746];
				12'd3747	: data <= weights[3747];
				12'd3748	: data <= weights[3748];
				12'd3749	: data <= weights[3749];
				12'd3750	: data <= weights[3750];
				12'd3751	: data <= weights[3751];
				12'd3752	: data <= weights[3752];
				12'd3753	: data <= weights[3753];
				12'd3754	: data <= weights[3754];
				12'd3755	: data <= weights[3755];
				12'd3756	: data <= weights[3756];
				12'd3757	: data <= weights[3757];
				12'd3758	: data <= weights[3758];
				12'd3759	: data <= weights[3759];
				12'd3760	: data <= weights[3760];
				12'd3761	: data <= weights[3761];
				12'd3762	: data <= weights[3762];
				12'd3763	: data <= weights[3763];
				12'd3764	: data <= weights[3764];
				12'd3765	: data <= weights[3765];
				12'd3766	: data <= weights[3766];
				12'd3767	: data <= weights[3767];
				12'd3768	: data <= weights[3768];
				12'd3769	: data <= weights[3769];
				12'd3770	: data <= weights[3770];
				12'd3771	: data <= weights[3771];
				12'd3772	: data <= weights[3772];
				12'd3773	: data <= weights[3773];
				12'd3774	: data <= weights[3774];
				12'd3775	: data <= weights[3775];
				12'd3776	: data <= weights[3776];
				12'd3777	: data <= weights[3777];
				12'd3778	: data <= weights[3778];
				12'd3779	: data <= weights[3779];
				12'd3780	: data <= weights[3780];
				12'd3781	: data <= weights[3781];
				12'd3782	: data <= weights[3782];
				12'd3783	: data <= weights[3783];
				12'd3784	: data <= weights[3784];
				12'd3785	: data <= weights[3785];
				12'd3786	: data <= weights[3786];
				12'd3787	: data <= weights[3787];
				12'd3788	: data <= weights[3788];
				12'd3789	: data <= weights[3789];
				12'd3790	: data <= weights[3790];
				12'd3791	: data <= weights[3791];
				12'd3792	: data <= weights[3792];
				12'd3793	: data <= weights[3793];
				12'd3794	: data <= weights[3794];
				12'd3795	: data <= weights[3795];
				12'd3796	: data <= weights[3796];
				12'd3797	: data <= weights[3797];
				12'd3798	: data <= weights[3798];
				12'd3799	: data <= weights[3799];
				12'd3800	: data <= weights[3800];
				12'd3801	: data <= weights[3801];
				12'd3802	: data <= weights[3802];
				12'd3803	: data <= weights[3803];
				12'd3804	: data <= weights[3804];
				12'd3805	: data <= weights[3805];
				12'd3806	: data <= weights[3806];
				12'd3807	: data <= weights[3807];
				12'd3808	: data <= weights[3808];
				12'd3809	: data <= weights[3809];
				12'd3810	: data <= weights[3810];
				12'd3811	: data <= weights[3811];
				12'd3812	: data <= weights[3812];
				12'd3813	: data <= weights[3813];
				12'd3814	: data <= weights[3814];
				12'd3815	: data <= weights[3815];
				12'd3816	: data <= weights[3816];
				12'd3817	: data <= weights[3817];
				12'd3818	: data <= weights[3818];
				12'd3819	: data <= weights[3819];
				12'd3820	: data <= weights[3820];
				12'd3821	: data <= weights[3821];
				12'd3822	: data <= weights[3822];
				12'd3823	: data <= weights[3823];
				12'd3824	: data <= weights[3824];
				12'd3825	: data <= weights[3825];
				12'd3826	: data <= weights[3826];
				12'd3827	: data <= weights[3827];
				12'd3828	: data <= weights[3828];
				12'd3829	: data <= weights[3829];
				12'd3830	: data <= weights[3830];
				12'd3831	: data <= weights[3831];
				12'd3832	: data <= weights[3832];
				12'd3833	: data <= weights[3833];
				12'd3834	: data <= weights[3834];
				12'd3835	: data <= weights[3835];
				12'd3836	: data <= weights[3836];
				12'd3837	: data <= weights[3837];
				12'd3838	: data <= weights[3838];
				12'd3839	: data <= weights[3839];
				12'd3840	: data <= weights[3840];
				12'd3841	: data <= weights[3841];
				12'd3842	: data <= weights[3842];
				12'd3843	: data <= weights[3843];
				12'd3844	: data <= weights[3844];
				12'd3845	: data <= weights[3845];
				12'd3846	: data <= weights[3846];
				12'd3847	: data <= weights[3847];
				12'd3848	: data <= weights[3848];
				12'd3849	: data <= weights[3849];
				12'd3850	: data <= weights[3850];
				12'd3851	: data <= weights[3851];
				12'd3852	: data <= weights[3852];
				12'd3853	: data <= weights[3853];
				12'd3854	: data <= weights[3854];
				12'd3855	: data <= weights[3855];
				12'd3856	: data <= weights[3856];
				12'd3857	: data <= weights[3857];
				12'd3858	: data <= weights[3858];
				12'd3859	: data <= weights[3859];
				12'd3860	: data <= weights[3860];
				12'd3861	: data <= weights[3861];
				12'd3862	: data <= weights[3862];
				12'd3863	: data <= weights[3863];
				12'd3864	: data <= weights[3864];
				12'd3865	: data <= weights[3865];
				12'd3866	: data <= weights[3866];
				12'd3867	: data <= weights[3867];
				12'd3868	: data <= weights[3868];
				12'd3869	: data <= weights[3869];
				12'd3870	: data <= weights[3870];
				12'd3871	: data <= weights[3871];
				12'd3872	: data <= weights[3872];
				12'd3873	: data <= weights[3873];
				12'd3874	: data <= weights[3874];
				12'd3875	: data <= weights[3875];
				12'd3876	: data <= weights[3876];
				12'd3877	: data <= weights[3877];
				12'd3878	: data <= weights[3878];
				12'd3879	: data <= weights[3879];
				12'd3880	: data <= weights[3880];
				12'd3881	: data <= weights[3881];
				12'd3882	: data <= weights[3882];
				12'd3883	: data <= weights[3883];
				12'd3884	: data <= weights[3884];
				12'd3885	: data <= weights[3885];
				12'd3886	: data <= weights[3886];
				12'd3887	: data <= weights[3887];
				12'd3888	: data <= weights[3888];
				12'd3889	: data <= weights[3889];
				12'd3890	: data <= weights[3890];
				12'd3891	: data <= weights[3891];
				12'd3892	: data <= weights[3892];
				12'd3893	: data <= weights[3893];
				12'd3894	: data <= weights[3894];
				12'd3895	: data <= weights[3895];
				12'd3896	: data <= weights[3896];
				12'd3897	: data <= weights[3897];
				12'd3898	: data <= weights[3898];
				12'd3899	: data <= weights[3899];
				12'd3900	: data <= weights[3900];
				12'd3901	: data <= weights[3901];
				12'd3902	: data <= weights[3902];
				12'd3903	: data <= weights[3903];
				12'd3904	: data <= weights[3904];
				12'd3905	: data <= weights[3905];
				12'd3906	: data <= weights[3906];
				12'd3907	: data <= weights[3907];
				12'd3908	: data <= weights[3908];
				12'd3909	: data <= weights[3909];
				12'd3910	: data <= weights[3910];
				12'd3911	: data <= weights[3911];
				12'd3912	: data <= weights[3912];
				12'd3913	: data <= weights[3913];
				12'd3914	: data <= weights[3914];
				12'd3915	: data <= weights[3915];
				12'd3916	: data <= weights[3916];
				12'd3917	: data <= weights[3917];
				12'd3918	: data <= weights[3918];
				12'd3919	: data <= weights[3919];
				12'd3920	: data <= weights[3920];
				12'd3921	: data <= weights[3921];
				12'd3922	: data <= weights[3922];
				12'd3923	: data <= weights[3923];
				12'd3924	: data <= weights[3924];
				12'd3925	: data <= weights[3925];
				12'd3926	: data <= weights[3926];
				12'd3927	: data <= weights[3927];
				12'd3928	: data <= weights[3928];
				12'd3929	: data <= weights[3929];
				12'd3930	: data <= weights[3930];
				12'd3931	: data <= weights[3931];
				12'd3932	: data <= weights[3932];
				12'd3933	: data <= weights[3933];
				12'd3934	: data <= weights[3934];
				12'd3935	: data <= weights[3935];
				12'd3936	: data <= weights[3936];
				12'd3937	: data <= weights[3937];
				12'd3938	: data <= weights[3938];
				12'd3939	: data <= weights[3939];
				12'd3940	: data <= weights[3940];
				12'd3941	: data <= weights[3941];
				12'd3942	: data <= weights[3942];
				12'd3943	: data <= weights[3943];
				12'd3944	: data <= weights[3944];
				12'd3945	: data <= weights[3945];
				12'd3946	: data <= weights[3946];
				12'd3947	: data <= weights[3947];
				12'd3948	: data <= weights[3948];
				12'd3949	: data <= weights[3949];
				12'd3950	: data <= weights[3950];
				12'd3951	: data <= weights[3951];
				12'd3952	: data <= weights[3952];
				12'd3953	: data <= weights[3953];
				12'd3954	: data <= weights[3954];
				12'd3955	: data <= weights[3955];
				12'd3956	: data <= weights[3956];
				12'd3957	: data <= weights[3957];
				12'd3958	: data <= weights[3958];
				12'd3959	: data <= weights[3959];
				12'd3960	: data <= weights[3960];
				12'd3961	: data <= weights[3961];
				12'd3962	: data <= weights[3962];
				12'd3963	: data <= weights[3963];
				12'd3964	: data <= weights[3964];
				12'd3965	: data <= weights[3965];
				12'd3966	: data <= weights[3966];
				12'd3967	: data <= weights[3967];
				12'd3968	: data <= weights[3968];
				12'd3969	: data <= weights[3969];
				12'd3970	: data <= weights[3970];
				12'd3971	: data <= weights[3971];
				12'd3972	: data <= weights[3972];
				12'd3973	: data <= weights[3973];
				12'd3974	: data <= weights[3974];
				12'd3975	: data <= weights[3975];
				12'd3976	: data <= weights[3976];
				12'd3977	: data <= weights[3977];
				12'd3978	: data <= weights[3978];
				12'd3979	: data <= weights[3979];
				12'd3980	: data <= weights[3980];
				12'd3981	: data <= weights[3981];
				12'd3982	: data <= weights[3982];
				12'd3983	: data <= weights[3983];
				12'd3984	: data <= weights[3984];
				12'd3985	: data <= weights[3985];
				12'd3986	: data <= weights[3986];
				12'd3987	: data <= weights[3987];
				12'd3988	: data <= weights[3988];
				12'd3989	: data <= weights[3989];
				12'd3990	: data <= weights[3990];
				12'd3991	: data <= weights[3991];
				12'd3992	: data <= weights[3992];
				12'd3993	: data <= weights[3993];
				12'd3994	: data <= weights[3994];
				12'd3995	: data <= weights[3995];
				12'd3996	: data <= weights[3996];
				12'd3997	: data <= weights[3997];
				12'd3998	: data <= weights[3998];
				12'd3999	: data <= weights[3999];
				12'd4000	: data <= weights[4000];
				12'd4001	: data <= weights[4001];
				12'd4002	: data <= weights[4002];
				12'd4003	: data <= weights[4003];
				12'd4004	: data <= weights[4004];
				12'd4005	: data <= weights[4005];
				12'd4006	: data <= weights[4006];
				12'd4007	: data <= weights[4007];
				12'd4008	: data <= weights[4008];
				12'd4009	: data <= weights[4009];
				12'd4010	: data <= weights[4010];
				12'd4011	: data <= weights[4011];
				12'd4012	: data <= weights[4012];
				12'd4013	: data <= weights[4013];
				12'd4014	: data <= weights[4014];
				12'd4015	: data <= weights[4015];
				12'd4016	: data <= weights[4016];
				12'd4017	: data <= weights[4017];
				12'd4018	: data <= weights[4018];
				12'd4019	: data <= weights[4019];
				12'd4020	: data <= weights[4020];
				12'd4021	: data <= weights[4021];
				12'd4022	: data <= weights[4022];
				12'd4023	: data <= weights[4023];
				12'd4024	: data <= weights[4024];
				12'd4025	: data <= weights[4025];
				12'd4026	: data <= weights[4026];
				12'd4027	: data <= weights[4027];
				12'd4028	: data <= weights[4028];
				12'd4029	: data <= weights[4029];
				12'd4030	: data <= weights[4030];
				12'd4031	: data <= weights[4031];
				12'd4032	: data <= weights[4032];
				12'd4033	: data <= weights[4033];
				12'd4034	: data <= weights[4034];
				12'd4035	: data <= weights[4035];
				12'd4036	: data <= weights[4036];
				12'd4037	: data <= weights[4037];
				12'd4038	: data <= weights[4038];
				12'd4039	: data <= weights[4039];
				12'd4040	: data <= weights[4040];
				12'd4041	: data <= weights[4041];
				12'd4042	: data <= weights[4042];
				12'd4043	: data <= weights[4043];
				12'd4044	: data <= weights[4044];
				12'd4045	: data <= weights[4045];
				12'd4046	: data <= weights[4046];
				12'd4047	: data <= weights[4047];
				12'd4048	: data <= weights[4048];
				12'd4049	: data <= weights[4049];
				12'd4050	: data <= weights[4050];
				12'd4051	: data <= weights[4051];
				12'd4052	: data <= weights[4052];
				12'd4053	: data <= weights[4053];
				12'd4054	: data <= weights[4054];
				12'd4055	: data <= weights[4055];
				12'd4056	: data <= weights[4056];
				12'd4057	: data <= weights[4057];
				12'd4058	: data <= weights[4058];
				12'd4059	: data <= weights[4059];
				12'd4060	: data <= weights[4060];
				12'd4061	: data <= weights[4061];
				12'd4062	: data <= weights[4062];
				12'd4063	: data <= weights[4063];
				12'd4064	: data <= weights[4064];
				default		: data <= 16'd0;
			endcase
		end else begin
			data <= data;
		end
	end

endmodule