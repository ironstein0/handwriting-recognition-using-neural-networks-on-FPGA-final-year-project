module traffic_generator(
	input wire clk,
	input wire [7:0] input_data