module ROM(
	input wire clk,
	input wire enable,
	input wire [11:0] address,
	output reg [15:0] data1,
	output reg [15:0] data2
	);

	reg [15:0] weights [4050:0];

	initial begin
		weights[0] <= 184;
		weights[1] <= 218;
		weights[2] <= 195;
		weights[3] <= 107;
		weights[4] <= 131;
		weights[5] <= 237;
		weights[6] <= 76;
		weights[7] <= 238;
		weights[8] <= 205;
		weights[9] <= 68;
		weights[10] <= 88;
		weights[11] <= 55;
		weights[12] <= 102;
		weights[13] <= 108;
		weights[14] <= 65;
		weights[15] <= 170;
		weights[16] <= 119;
		weights[17] <= 125;
		weights[18] <= 79;
		weights[19] <= 231;
		weights[20] <= 203;
		weights[21] <= 5;
		weights[22] <= 100;
		weights[23] <= 213;
		weights[24] <= 124;
		weights[25] <= 56;
		weights[26] <= 166;
		weights[27] <= 35;
		weights[28] <= 139;
		weights[29] <= 135;
		weights[30] <= 225;
		weights[31] <= 119;
		weights[32] <= 170;
		weights[33] <= 193;
		weights[34] <= 125;
		weights[35] <= 227;
		weights[36] <= 116;
		weights[37] <= 159;
		weights[38] <= 230;
		weights[39] <= 128;
		weights[40] <= 192;
		weights[41] <= 25;
		weights[42] <= 187;
		weights[43] <= 80;
		weights[44] <= 116;
		weights[45] <= 133;
		weights[46] <= 103;
		weights[47] <= 229;
		weights[48] <= 147;
		weights[49] <= 201;
		weights[50] <= 177;
		weights[51] <= 161;
		weights[52] <= 135;
		weights[53] <= 146;
		weights[54] <= 1;
		weights[55] <= 228;
		weights[56] <= 239;
		weights[57] <= 54;
		weights[58] <= 82;
		weights[59] <= 12;
		weights[60] <= 51;
		weights[61] <= 142;
		weights[62] <= 52;
		weights[63] <= 172;
		weights[64] <= 129;
		weights[65] <= 91;
		weights[66] <= 56;
		weights[67] <= 170;
		weights[68] <= 247;
		weights[69] <= 102;
		weights[70] <= 13;
		weights[71] <= 137;
		weights[72] <= 212;
		weights[73] <= 200;
		weights[74] <= 51;
		weights[75] <= 155;
		weights[76] <= 173;
		weights[77] <= 137;
		weights[78] <= 55;
		weights[79] <= 117;
		weights[80] <= 174;
		weights[81] <= 63;
		weights[82] <= 241;
		weights[83] <= 21;
		weights[84] <= 58;
		weights[85] <= 22;
		weights[86] <= 88;
		weights[87] <= 227;
		weights[88] <= 94;
		weights[89] <= 194;
		weights[90] <= 118;
		weights[91] <= 22;
		weights[92] <= 172;
		weights[93] <= 232;
		weights[94] <= 247;
		weights[95] <= 45;
		weights[96] <= 88;
		weights[97] <= 143;
		weights[98] <= 51;
		weights[99] <= 106;
		weights[100] <= 212;
		weights[101] <= 244;
		weights[102] <= 246;
		weights[103] <= 245;
		weights[104] <= 166;
		weights[105] <= 157;
		weights[106] <= 143;
		weights[107] <= 249;
		weights[108] <= 111;
		weights[109] <= 30;
		weights[110] <= 110;
		weights[111] <= 168;
		weights[112] <= 117;
		weights[113] <= 13;
		weights[114] <= 58;
		weights[115] <= 140;
		weights[116] <= 255;
		weights[117] <= 170;
		weights[118] <= 136;
		weights[119] <= 214;
		weights[120] <= 91;
		weights[121] <= 27;
		weights[122] <= 142;
		weights[123] <= 126;
		weights[124] <= 228;
		weights[125] <= 54;
		weights[126] <= 176;
		weights[127] <= 139;
		weights[128] <= 187;
		weights[129] <= 150;
		weights[130] <= 16;
		weights[131] <= 62;
		weights[132] <= 44;
		weights[133] <= 58;
		weights[134] <= 166;
		weights[135] <= 168;
		weights[136] <= 151;
		weights[137] <= 1;
		weights[138] <= 56;
		weights[139] <= 50;
		weights[140] <= 41;
		weights[141] <= 187;
		weights[142] <= 142;
		weights[143] <= 151;
		weights[144] <= 190;
		weights[145] <= 15;
		weights[146] <= 171;
		weights[147] <= 54;
		weights[148] <= 33;
		weights[149] <= 146;
		weights[150] <= 40;
		weights[151] <= 69;
		weights[152] <= 36;
		weights[153] <= 100;
		weights[154] <= 30;
		weights[155] <= 246;
		weights[156] <= 171;
		weights[157] <= 207;
		weights[158] <= 162;
		weights[159] <= 85;
		weights[160] <= 57;
		weights[161] <= 22;
		weights[162] <= 53;
		weights[163] <= 155;
		weights[164] <= 63;
		weights[165] <= 246;
		weights[166] <= 48;
		weights[167] <= 64;
		weights[168] <= 70;
		weights[169] <= 191;
		weights[170] <= 88;
		weights[171] <= 119;
		weights[172] <= 75;
		weights[173] <= 67;
		weights[174] <= 197;
		weights[175] <= 110;
		weights[176] <= 7;
		weights[177] <= 168;
		weights[178] <= 217;
		weights[179] <= 35;
		weights[180] <= 162;
		weights[181] <= 25;
		weights[182] <= 189;
		weights[183] <= 222;
		weights[184] <= 29;
		weights[185] <= 199;
		weights[186] <= 200;
		weights[187] <= 224;
		weights[188] <= 29;
		weights[189] <= 250;
		weights[190] <= 82;
		weights[191] <= 145;
		weights[192] <= 129;
		weights[193] <= 175;
		weights[194] <= 58;
		weights[195] <= 105;
		weights[196] <= 50;
		weights[197] <= 132;
		weights[198] <= 11;
		weights[199] <= 103;
		weights[200] <= 39;
		weights[201] <= 75;
		weights[202] <= 255;
		weights[203] <= 10;
		weights[204] <= 64;
		weights[205] <= 178;
		weights[206] <= 242;
		weights[207] <= 162;
		weights[208] <= 8;
		weights[209] <= 219;
		weights[210] <= 89;
		weights[211] <= 194;
		weights[212] <= 129;
		weights[213] <= 246;
		weights[214] <= 245;
		weights[215] <= 13;
		weights[216] <= 76;
		weights[217] <= 192;
		weights[218] <= 161;
		weights[219] <= 35;
		weights[220] <= 120;
		weights[221] <= 238;
		weights[222] <= 16;
		weights[223] <= 119;
		weights[224] <= 118;
		weights[225] <= 175;
		weights[226] <= 90;
		weights[227] <= 172;
		weights[228] <= 43;
		weights[229] <= 139;
		weights[230] <= 5;
		weights[231] <= 33;
		weights[232] <= 70;
		weights[233] <= 196;
		weights[234] <= 178;
		weights[235] <= 96;
		weights[236] <= 116;
		weights[237] <= 227;
		weights[238] <= 137;
		weights[239] <= 197;
		weights[240] <= 187;
		weights[241] <= 214;
		weights[242] <= 117;
		weights[243] <= 204;
		weights[244] <= 68;
		weights[245] <= 187;
		weights[246] <= 35;
		weights[247] <= 55;
		weights[248] <= 71;
		weights[249] <= 45;
		weights[250] <= 114;
		weights[251] <= 143;
		weights[252] <= 148;
		weights[253] <= 175;
		weights[254] <= 137;
		weights[255] <= 209;
		weights[256] <= 109;
		weights[257] <= 206;
		weights[258] <= 73;
		weights[259] <= 50;
		weights[260] <= 20;
		weights[261] <= 178;
		weights[262] <= 192;
		weights[263] <= 45;
		weights[264] <= 147;
		weights[265] <= 78;
		weights[266] <= 169;
		weights[267] <= 155;
		weights[268] <= 255;
		weights[269] <= 94;
		weights[270] <= 88;
		weights[271] <= 90;
		weights[272] <= 45;
		weights[273] <= 82;
		weights[274] <= 14;
		weights[275] <= 140;
		weights[276] <= 122;
		weights[277] <= 184;
		weights[278] <= 25;
		weights[279] <= 199;
		weights[280] <= 132;
		weights[281] <= 134;
		weights[282] <= 60;
		weights[283] <= 239;
		weights[284] <= 130;
		weights[285] <= 192;
		weights[286] <= 86;
		weights[287] <= 213;
		weights[288] <= 35;
		weights[289] <= 125;
		weights[290] <= 178;
		weights[291] <= 189;
		weights[292] <= 66;
		weights[293] <= 237;
		weights[294] <= 156;
		weights[295] <= 94;
		weights[296] <= 213;
		weights[297] <= 125;
		weights[298] <= 155;
		weights[299] <= 207;
		weights[300] <= 221;
		weights[301] <= 10;
		weights[302] <= 48;
		weights[303] <= 4;
		weights[304] <= 200;
		weights[305] <= 194;
		weights[306] <= 61;
		weights[307] <= 113;
		weights[308] <= 104;
		weights[309] <= 33;
		weights[310] <= 189;
		weights[311] <= 14;
		weights[312] <= 213;
		weights[313] <= 254;
		weights[314] <= 120;
		weights[315] <= 227;
		weights[316] <= 105;
		weights[317] <= 24;
		weights[318] <= 153;
		weights[319] <= 215;
		weights[320] <= 21;
		weights[321] <= 213;
		weights[322] <= 134;
		weights[323] <= 50;
		weights[324] <= 47;
		weights[325] <= 170;
		weights[326] <= 236;
		weights[327] <= 213;
		weights[328] <= 136;
		weights[329] <= 149;
		weights[330] <= 138;
		weights[331] <= 199;
		weights[332] <= 214;
		weights[333] <= 80;
		weights[334] <= 226;
		weights[335] <= 232;
		weights[336] <= 181;
		weights[337] <= 18;
		weights[338] <= 65;
		weights[339] <= 140;
		weights[340] <= 215;
		weights[341] <= 16;
		weights[342] <= 26;
		weights[343] <= 71;
		weights[344] <= 26;
		weights[345] <= 76;
		weights[346] <= 121;
		weights[347] <= 105;
		weights[348] <= 209;
		weights[349] <= 180;
		weights[350] <= 92;
		weights[351] <= 141;
		weights[352] <= 154;
		weights[353] <= 196;
		weights[354] <= 99;
		weights[355] <= 60;
		weights[356] <= 179;
		weights[357] <= 195;
		weights[358] <= 6;
		weights[359] <= 17;
		weights[360] <= 55;
		weights[361] <= 254;
		weights[362] <= 222;
		weights[363] <= 18;
		weights[364] <= 210;
		weights[365] <= 105;
		weights[366] <= 54;
		weights[367] <= 131;
		weights[368] <= 143;
		weights[369] <= 237;
		weights[370] <= 239;
		weights[371] <= 153;
		weights[372] <= 88;
		weights[373] <= 110;
		weights[374] <= 197;
		weights[375] <= 24;
		weights[376] <= 124;
		weights[377] <= 40;
		weights[378] <= 117;
		weights[379] <= 52;
		weights[380] <= 211;
		weights[381] <= 41;
		weights[382] <= 15;
		weights[383] <= 154;
		weights[384] <= 225;
		weights[385] <= 182;
		weights[386] <= 118;
		weights[387] <= 241;
		weights[388] <= 161;
		weights[389] <= 237;
		weights[390] <= 230;
		weights[391] <= 145;
		weights[392] <= 213;
		weights[393] <= 200;
		weights[394] <= 121;
		weights[395] <= 107;
		weights[396] <= 77;
		weights[397] <= 46;
		weights[398] <= 80;
		weights[399] <= 4;
		weights[400] <= 102;
		weights[401] <= 155;
		weights[402] <= 180;
		weights[403] <= 112;
		weights[404] <= 186;
		weights[405] <= 107;
		weights[406] <= 46;
		weights[407] <= 127;
		weights[408] <= 33;
		weights[409] <= 193;
		weights[410] <= 180;
		weights[411] <= 139;
		weights[412] <= 36;
		weights[413] <= 4;
		weights[414] <= 131;
		weights[415] <= 249;
		weights[416] <= 158;
		weights[417] <= 64;
		weights[418] <= 12;
		weights[419] <= 21;
		weights[420] <= 69;
		weights[421] <= 69;
		weights[422] <= 110;
		weights[423] <= 27;
		weights[424] <= 192;
		weights[425] <= 246;
		weights[426] <= 152;
		weights[427] <= 49;
		weights[428] <= 147;
		weights[429] <= 64;
		weights[430] <= 188;
		weights[431] <= 154;
		weights[432] <= 196;
		weights[433] <= 254;
		weights[434] <= 24;
		weights[435] <= 41;
		weights[436] <= 153;
		weights[437] <= 86;
		weights[438] <= 58;
		weights[439] <= 69;
		weights[440] <= 108;
		weights[441] <= 106;
		weights[442] <= 164;
		weights[443] <= 202;
		weights[444] <= 41;
		weights[445] <= 73;
		weights[446] <= 219;
		weights[447] <= 182;
		weights[448] <= 54;
		weights[449] <= 103;
		weights[450] <= 150;
		weights[451] <= 65;
		weights[452] <= 134;
		weights[453] <= 12;
		weights[454] <= 130;
		weights[455] <= 131;
		weights[456] <= 239;
		weights[457] <= 224;
		weights[458] <= 49;
		weights[459] <= 242;
		weights[460] <= 38;
		weights[461] <= 200;
		weights[462] <= 216;
		weights[463] <= 184;
		weights[464] <= 186;
		weights[465] <= 230;
		weights[466] <= 8;
		weights[467] <= 150;
		weights[468] <= 107;
		weights[469] <= 174;
		weights[470] <= 9;
		weights[471] <= 54;
		weights[472] <= 164;
		weights[473] <= 244;
		weights[474] <= 20;
		weights[475] <= 116;
		weights[476] <= 216;
		weights[477] <= 84;
		weights[478] <= 236;
		weights[479] <= 112;
		weights[480] <= 86;
		weights[481] <= 124;
		weights[482] <= 120;
		weights[483] <= 112;
		weights[484] <= 223;
		weights[485] <= 31;
		weights[486] <= 195;
		weights[487] <= 13;
		weights[488] <= 238;
		weights[489] <= 114;
		weights[490] <= 114;
		weights[491] <= 13;
		weights[492] <= 214;
		weights[493] <= 46;
		weights[494] <= 233;
		weights[495] <= 194;
		weights[496] <= 52;
		weights[497] <= 170;
		weights[498] <= 191;
		weights[499] <= 173;
		weights[500] <= 134;
		weights[501] <= 236;
		weights[502] <= 105;
		weights[503] <= 86;
		weights[504] <= 167;
		weights[505] <= 181;
		weights[506] <= 150;
		weights[507] <= 156;
		weights[508] <= 49;
		weights[509] <= 142;
		weights[510] <= 156;
		weights[511] <= 254;
		weights[512] <= 18;
		weights[513] <= 57;
		weights[514] <= 141;
		weights[515] <= 26;
		weights[516] <= 22;
		weights[517] <= 184;
		weights[518] <= 65;
		weights[519] <= 14;
		weights[520] <= 171;
		weights[521] <= 160;
		weights[522] <= 112;
		weights[523] <= 101;
		weights[524] <= 248;
		weights[525] <= 1;
		weights[526] <= 175;
		weights[527] <= 14;
		weights[528] <= 199;
		weights[529] <= 27;
		weights[530] <= 213;
		weights[531] <= 61;
		weights[532] <= 232;
		weights[533] <= 245;
		weights[534] <= 195;
		weights[535] <= 89;
		weights[536] <= 33;
		weights[537] <= 12;
		weights[538] <= 187;
		weights[539] <= 121;
		weights[540] <= 85;
		weights[541] <= 191;
		weights[542] <= 91;
		weights[543] <= 235;
		weights[544] <= 209;
		weights[545] <= 224;
		weights[546] <= 102;
		weights[547] <= 31;
		weights[548] <= 176;
		weights[549] <= 235;
		weights[550] <= 192;
		weights[551] <= 152;
		weights[552] <= 138;
		weights[553] <= 165;
		weights[554] <= 138;
		weights[555] <= 223;
		weights[556] <= 190;
		weights[557] <= 25;
		weights[558] <= 111;
		weights[559] <= 234;
		weights[560] <= 206;
		weights[561] <= 33;
		weights[562] <= 161;
		weights[563] <= 215;
		weights[564] <= 229;
		weights[565] <= 180;
		weights[566] <= 1;
		weights[567] <= 182;
		weights[568] <= 92;
		weights[569] <= 237;
		weights[570] <= 136;
		weights[571] <= 64;
		weights[572] <= 122;
		weights[573] <= 247;
		weights[574] <= 121;
		weights[575] <= 132;
		weights[576] <= 106;
		weights[577] <= 18;
		weights[578] <= 227;
		weights[579] <= 115;
		weights[580] <= 25;
		weights[581] <= 207;
		weights[582] <= 186;
		weights[583] <= 39;
		weights[584] <= 32;
		weights[585] <= 174;
		weights[586] <= 31;
		weights[587] <= 226;
		weights[588] <= 173;
		weights[589] <= 117;
		weights[590] <= 92;
		weights[591] <= 208;
		weights[592] <= 19;
		weights[593] <= 188;
		weights[594] <= 60;
		weights[595] <= 74;
		weights[596] <= 248;
		weights[597] <= 105;
		weights[598] <= 143;
		weights[599] <= 47;
		weights[600] <= 25;
		weights[601] <= 227;
		weights[602] <= 209;
		weights[603] <= 219;
		weights[604] <= 89;
		weights[605] <= 208;
		weights[606] <= 38;
		weights[607] <= 8;
		weights[608] <= 106;
		weights[609] <= 93;
		weights[610] <= 230;
		weights[611] <= 34;
		weights[612] <= 193;
		weights[613] <= 161;
		weights[614] <= 30;
		weights[615] <= 151;
		weights[616] <= 119;
		weights[617] <= 89;
		weights[618] <= 185;
		weights[619] <= 15;
		weights[620] <= 158;
		weights[621] <= 231;
		weights[622] <= 242;
		weights[623] <= 255;
		weights[624] <= 229;
		weights[625] <= 93;
		weights[626] <= 166;
		weights[627] <= 215;
		weights[628] <= 85;
		weights[629] <= 2;
		weights[630] <= 171;
		weights[631] <= 53;
		weights[632] <= 84;
		weights[633] <= 209;
		weights[634] <= 141;
		weights[635] <= 46;
		weights[636] <= 128;
		weights[637] <= 72;
		weights[638] <= 190;
		weights[639] <= 76;
		weights[640] <= 95;
		weights[641] <= 38;
		weights[642] <= 225;
		weights[643] <= 204;
		weights[644] <= 1;
		weights[645] <= 50;
		weights[646] <= 76;
		weights[647] <= 96;
		weights[648] <= 88;
		weights[649] <= 55;
		weights[650] <= 77;
		weights[651] <= 150;
		weights[652] <= 150;
		weights[653] <= 32;
		weights[654] <= 189;
		weights[655] <= 24;
		weights[656] <= 151;
		weights[657] <= 13;
		weights[658] <= 254;
		weights[659] <= 38;
		weights[660] <= 199;
		weights[661] <= 80;
		weights[662] <= 241;
		weights[663] <= 133;
		weights[664] <= 76;
		weights[665] <= 94;
		weights[666] <= 125;
		weights[667] <= 98;
		weights[668] <= 229;
		weights[669] <= 96;
		weights[670] <= 215;
		weights[671] <= 191;
		weights[672] <= 62;
		weights[673] <= 248;
		weights[674] <= 210;
		weights[675] <= 138;
		weights[676] <= 109;
		weights[677] <= 59;
		weights[678] <= 156;
		weights[679] <= 99;
		weights[680] <= 128;
		weights[681] <= 156;
		weights[682] <= 70;
		weights[683] <= 202;
		weights[684] <= 32;
		weights[685] <= 186;
		weights[686] <= 78;
		weights[687] <= 231;
		weights[688] <= 251;
		weights[689] <= 99;
		weights[690] <= 189;
		weights[691] <= 132;
		weights[692] <= 114;
		weights[693] <= 39;
		weights[694] <= 213;
		weights[695] <= 232;
		weights[696] <= 206;
		weights[697] <= 104;
		weights[698] <= 133;
		weights[699] <= 255;
		weights[700] <= 26;
		weights[701] <= 163;
		weights[702] <= 195;
		weights[703] <= 191;
		weights[704] <= 101;
		weights[705] <= 41;
		weights[706] <= 251;
		weights[707] <= 252;
		weights[708] <= 117;
		weights[709] <= 16;
		weights[710] <= 100;
		weights[711] <= 42;
		weights[712] <= 8;
		weights[713] <= 152;
		weights[714] <= 153;
		weights[715] <= 113;
		weights[716] <= 206;
		weights[717] <= 67;
		weights[718] <= 14;
		weights[719] <= 160;
		weights[720] <= 64;
		weights[721] <= 221;
		weights[722] <= 88;
		weights[723] <= 104;
		weights[724] <= 68;
		weights[725] <= 255;
		weights[726] <= 9;
		weights[727] <= 88;
		weights[728] <= 116;
		weights[729] <= 41;
		weights[730] <= 127;
		weights[731] <= 161;
		weights[732] <= 124;
		weights[733] <= 16;
		weights[734] <= 148;
		weights[735] <= 66;
		weights[736] <= 93;
		weights[737] <= 3;
		weights[738] <= 205;
		weights[739] <= 85;
		weights[740] <= 73;
		weights[741] <= 135;
		weights[742] <= 114;
		weights[743] <= 108;
		weights[744] <= 229;
		weights[745] <= 173;
		weights[746] <= 13;
		weights[747] <= 141;
		weights[748] <= 46;
		weights[749] <= 91;
		weights[750] <= 189;
		weights[751] <= 119;
		weights[752] <= 47;
		weights[753] <= 76;
		weights[754] <= 195;
		weights[755] <= 194;
		weights[756] <= 191;
		weights[757] <= 83;
		weights[758] <= 27;
		weights[759] <= 120;
		weights[760] <= 11;
		weights[761] <= 41;
		weights[762] <= 161;
		weights[763] <= 64;
		weights[764] <= 41;
		weights[765] <= 149;
		weights[766] <= 189;
		weights[767] <= 24;
		weights[768] <= 156;
		weights[769] <= 125;
		weights[770] <= 36;
		weights[771] <= 251;
		weights[772] <= 130;
		weights[773] <= 52;
		weights[774] <= 12;
		weights[775] <= 170;
		weights[776] <= 59;
		weights[777] <= 183;
		weights[778] <= 118;
		weights[779] <= 127;
		weights[780] <= 71;
		weights[781] <= 47;
		weights[782] <= 126;
		weights[783] <= 216;
		weights[784] <= 123;
		weights[785] <= 44;
		weights[786] <= 209;
		weights[787] <= 70;
		weights[788] <= 189;
		weights[789] <= 22;
		weights[790] <= 71;
		weights[791] <= 155;
		weights[792] <= 9;
		weights[793] <= 252;
		weights[794] <= 232;
		weights[795] <= 83;
		weights[796] <= 24;
		weights[797] <= 123;
		weights[798] <= 117;
		weights[799] <= 108;
		weights[800] <= 204;
		weights[801] <= 34;
		weights[802] <= 96;
		weights[803] <= 24;
		weights[804] <= 56;
		weights[805] <= 72;
		weights[806] <= 228;
		weights[807] <= 78;
		weights[808] <= 221;
		weights[809] <= 45;
		weights[810] <= 254;
		weights[811] <= 36;
		weights[812] <= 51;
		weights[813] <= 208;
		weights[814] <= 18;
		weights[815] <= 164;
		weights[816] <= 91;
		weights[817] <= 232;
		weights[818] <= 1;
		weights[819] <= 254;
		weights[820] <= 55;
		weights[821] <= 210;
		weights[822] <= 219;
		weights[823] <= 220;
		weights[824] <= 154;
		weights[825] <= 6;
		weights[826] <= 69;
		weights[827] <= 43;
		weights[828] <= 139;
		weights[829] <= 248;
		weights[830] <= 56;
		weights[831] <= 126;
		weights[832] <= 153;
		weights[833] <= 213;
		weights[834] <= 96;
		weights[835] <= 7;
		weights[836] <= 22;
		weights[837] <= 174;
		weights[838] <= 162;
		weights[839] <= 96;
		weights[840] <= 240;
		weights[841] <= 149;
		weights[842] <= 30;
		weights[843] <= 157;
		weights[844] <= 37;
		weights[845] <= 174;
		weights[846] <= 156;
		weights[847] <= 136;
		weights[848] <= 225;
		weights[849] <= 122;
		weights[850] <= 5;
		weights[851] <= 203;
		weights[852] <= 51;
		weights[853] <= 215;
		weights[854] <= 22;
		weights[855] <= 160;
		weights[856] <= 199;
		weights[857] <= 111;
		weights[858] <= 118;
		weights[859] <= 104;
		weights[860] <= 221;
		weights[861] <= 101;
		weights[862] <= 145;
		weights[863] <= 166;
		weights[864] <= 166;
		weights[865] <= 167;
		weights[866] <= 44;
		weights[867] <= 52;
		weights[868] <= 175;
		weights[869] <= 178;
		weights[870] <= 222;
		weights[871] <= 112;
		weights[872] <= 243;
		weights[873] <= 94;
		weights[874] <= 83;
		weights[875] <= 100;
		weights[876] <= 214;
		weights[877] <= 234;
		weights[878] <= 175;
		weights[879] <= 32;
		weights[880] <= 249;
		weights[881] <= 62;
		weights[882] <= 193;
		weights[883] <= 190;
		weights[884] <= 125;
		weights[885] <= 96;
		weights[886] <= 222;
		weights[887] <= 41;
		weights[888] <= 124;
		weights[889] <= 20;
		weights[890] <= 32;
		weights[891] <= 132;
		weights[892] <= 91;
		weights[893] <= 41;
		weights[894] <= 243;
		weights[895] <= 250;
		weights[896] <= 233;
		weights[897] <= 106;
		weights[898] <= 101;
		weights[899] <= 86;
		weights[900] <= 145;
		weights[901] <= 187;
		weights[902] <= 239;
		weights[903] <= 240;
		weights[904] <= 112;
		weights[905] <= 3;
		weights[906] <= 239;
		weights[907] <= 63;
		weights[908] <= 32;
		weights[909] <= 150;
		weights[910] <= 102;
		weights[911] <= 4;
		weights[912] <= 224;
		weights[913] <= 78;
		weights[914] <= 213;
		weights[915] <= 61;
		weights[916] <= 149;
		weights[917] <= 50;
		weights[918] <= 211;
		weights[919] <= 247;
		weights[920] <= 156;
		weights[921] <= 191;
		weights[922] <= 236;
		weights[923] <= 244;
		weights[924] <= 108;
		weights[925] <= 191;
		weights[926] <= 115;
		weights[927] <= 128;
		weights[928] <= 76;
		weights[929] <= 99;
		weights[930] <= 99;
		weights[931] <= 218;
		weights[932] <= 184;
		weights[933] <= 60;
		weights[934] <= 59;
		weights[935] <= 5;
		weights[936] <= 145;
		weights[937] <= 148;
		weights[938] <= 193;
		weights[939] <= 188;
		weights[940] <= 26;
		weights[941] <= 208;
		weights[942] <= 129;
		weights[943] <= 203;
		weights[944] <= 208;
		weights[945] <= 159;
		weights[946] <= 227;
		weights[947] <= 134;
		weights[948] <= 11;
		weights[949] <= 8;
		weights[950] <= 190;
		weights[951] <= 220;
		weights[952] <= 77;
		weights[953] <= 247;
		weights[954] <= 105;
		weights[955] <= 115;
		weights[956] <= 127;
		weights[957] <= 143;
		weights[958] <= 180;
		weights[959] <= 122;
		weights[960] <= 154;
		weights[961] <= 66;
		weights[962] <= 229;
		weights[963] <= 127;
		weights[964] <= 40;
		weights[965] <= 17;
		weights[966] <= 74;
		weights[967] <= 255;
		weights[968] <= 87;
		weights[969] <= 206;
		weights[970] <= 162;
		weights[971] <= 123;
		weights[972] <= 185;
		weights[973] <= 154;
		weights[974] <= 41;
		weights[975] <= 188;
		weights[976] <= 244;
		weights[977] <= 81;
		weights[978] <= 96;
		weights[979] <= 146;
		weights[980] <= 132;
		weights[981] <= 169;
		weights[982] <= 105;
		weights[983] <= 89;
		weights[984] <= 87;
		weights[985] <= 208;
		weights[986] <= 77;
		weights[987] <= 206;
		weights[988] <= 231;
		weights[989] <= 71;
		weights[990] <= 50;
		weights[991] <= 46;
		weights[992] <= 105;
		weights[993] <= 239;
		weights[994] <= 248;
		weights[995] <= 108;
		weights[996] <= 80;
		weights[997] <= 185;
		weights[998] <= 179;
		weights[999] <= 193;
		weights[1000] <= 86;
		weights[1001] <= 210;
		weights[1002] <= 171;
		weights[1003] <= 134;
		weights[1004] <= 53;
		weights[1005] <= 84;
		weights[1006] <= 201;
		weights[1007] <= 12;
		weights[1008] <= 160;
		weights[1009] <= 22;
		weights[1010] <= 142;
		weights[1011] <= 208;
		weights[1012] <= 77;
		weights[1013] <= 79;
		weights[1014] <= 122;
		weights[1015] <= 137;
		weights[1016] <= 29;
		weights[1017] <= 229;
		weights[1018] <= 133;
		weights[1019] <= 65;
		weights[1020] <= 35;
		weights[1021] <= 11;
		weights[1022] <= 20;
		weights[1023] <= 165;
		weights[1024] <= 82;
		weights[1025] <= 79;
		weights[1026] <= 34;
		weights[1027] <= 53;
		weights[1028] <= 40;
		weights[1029] <= 238;
		weights[1030] <= 110;
		weights[1031] <= 244;
		weights[1032] <= 249;
		weights[1033] <= 80;
		weights[1034] <= 146;
		weights[1035] <= 96;
		weights[1036] <= 86;
		weights[1037] <= 197;
		weights[1038] <= 32;
		weights[1039] <= 246;
		weights[1040] <= 165;
		weights[1041] <= 47;
		weights[1042] <= 83;
		weights[1043] <= 26;
		weights[1044] <= 227;
		weights[1045] <= 100;
		weights[1046] <= 117;
		weights[1047] <= 80;
		weights[1048] <= 115;
		weights[1049] <= 110;
		weights[1050] <= 30;
		weights[1051] <= 158;
		weights[1052] <= 86;
		weights[1053] <= 14;
		weights[1054] <= 172;
		weights[1055] <= 216;
		weights[1056] <= 245;
		weights[1057] <= 194;
		weights[1058] <= 246;
		weights[1059] <= 248;
		weights[1060] <= 156;
		weights[1061] <= 73;
		weights[1062] <= 94;
		weights[1063] <= 154;
		weights[1064] <= 227;
		weights[1065] <= 116;
		weights[1066] <= 184;
		weights[1067] <= 30;
		weights[1068] <= 186;
		weights[1069] <= 171;
		weights[1070] <= 180;
		weights[1071] <= 133;
		weights[1072] <= 10;
		weights[1073] <= 176;
		weights[1074] <= 146;
		weights[1075] <= 3;
		weights[1076] <= 210;
		weights[1077] <= 170;
		weights[1078] <= 229;
		weights[1079] <= 126;
		weights[1080] <= 155;
		weights[1081] <= 53;
		weights[1082] <= 32;
		weights[1083] <= 248;
		weights[1084] <= 89;
		weights[1085] <= 165;
		weights[1086] <= 141;
		weights[1087] <= 113;
		weights[1088] <= 206;
		weights[1089] <= 206;
		weights[1090] <= 25;
		weights[1091] <= 131;
		weights[1092] <= 227;
		weights[1093] <= 115;
		weights[1094] <= 51;
		weights[1095] <= 22;
		weights[1096] <= 192;
		weights[1097] <= 141;
		weights[1098] <= 158;
		weights[1099] <= 75;
		weights[1100] <= 137;
		weights[1101] <= 49;
		weights[1102] <= 151;
		weights[1103] <= 94;
		weights[1104] <= 87;
		weights[1105] <= 38;
		weights[1106] <= 132;
		weights[1107] <= 96;
		weights[1108] <= 144;
		weights[1109] <= 78;
		weights[1110] <= 247;
		weights[1111] <= 78;
		weights[1112] <= 242;
		weights[1113] <= 107;
		weights[1114] <= 104;
		weights[1115] <= 112;
		weights[1116] <= 1;
		weights[1117] <= 13;
		weights[1118] <= 94;
		weights[1119] <= 13;
		weights[1120] <= 175;
		weights[1121] <= 161;
		weights[1122] <= 100;
		weights[1123] <= 144;
		weights[1124] <= 32;
		weights[1125] <= 181;
		weights[1126] <= 149;
		weights[1127] <= 159;
		weights[1128] <= 187;
		weights[1129] <= 138;
		weights[1130] <= 182;
		weights[1131] <= 208;
		weights[1132] <= 109;
		weights[1133] <= 16;
		weights[1134] <= 26;
		weights[1135] <= 59;
		weights[1136] <= 1;
		weights[1137] <= 41;
		weights[1138] <= 93;
		weights[1139] <= 131;
		weights[1140] <= 18;
		weights[1141] <= 95;
		weights[1142] <= 130;
		weights[1143] <= 220;
		weights[1144] <= 17;
		weights[1145] <= 193;
		weights[1146] <= 146;
		weights[1147] <= 124;
		weights[1148] <= 112;
		weights[1149] <= 131;
		weights[1150] <= 47;
		weights[1151] <= 18;
		weights[1152] <= 47;
		weights[1153] <= 162;
		weights[1154] <= 214;
		weights[1155] <= 174;
		weights[1156] <= 73;
		weights[1157] <= 198;
		weights[1158] <= 244;
		weights[1159] <= 63;
		weights[1160] <= 6;
		weights[1161] <= 172;
		weights[1162] <= 26;
		weights[1163] <= 144;
		weights[1164] <= 97;
		weights[1165] <= 97;
		weights[1166] <= 66;
		weights[1167] <= 130;
		weights[1168] <= 116;
		weights[1169] <= 217;
		weights[1170] <= 66;
		weights[1171] <= 33;
		weights[1172] <= 99;
		weights[1173] <= 128;
		weights[1174] <= 83;
		weights[1175] <= 11;
		weights[1176] <= 148;
		weights[1177] <= 247;
		weights[1178] <= 216;
		weights[1179] <= 93;
		weights[1180] <= 108;
		weights[1181] <= 240;
		weights[1182] <= 203;
		weights[1183] <= 84;
		weights[1184] <= 140;
		weights[1185] <= 202;
		weights[1186] <= 85;
		weights[1187] <= 16;
		weights[1188] <= 80;
		weights[1189] <= 75;
		weights[1190] <= 230;
		weights[1191] <= 228;
		weights[1192] <= 144;
		weights[1193] <= 135;
		weights[1194] <= 235;
		weights[1195] <= 162;
		weights[1196] <= 79;
		weights[1197] <= 200;
		weights[1198] <= 100;
		weights[1199] <= 191;
		weights[1200] <= 80;
		weights[1201] <= 13;
		weights[1202] <= 60;
		weights[1203] <= 124;
		weights[1204] <= 163;
		weights[1205] <= 255;
		weights[1206] <= 119;
		weights[1207] <= 161;
		weights[1208] <= 132;
		weights[1209] <= 245;
		weights[1210] <= 14;
		weights[1211] <= 97;
		weights[1212] <= 254;
		weights[1213] <= 73;
		weights[1214] <= 82;
		weights[1215] <= 123;
		weights[1216] <= 60;
		weights[1217] <= 84;
		weights[1218] <= 122;
		weights[1219] <= 150;
		weights[1220] <= 225;
		weights[1221] <= 91;
		weights[1222] <= 47;
		weights[1223] <= 130;
		weights[1224] <= 239;
		weights[1225] <= 240;
		weights[1226] <= 112;
		weights[1227] <= 119;
		weights[1228] <= 61;
		weights[1229] <= 71;
		weights[1230] <= 148;
		weights[1231] <= 116;
		weights[1232] <= 234;
		weights[1233] <= 158;
		weights[1234] <= 165;
		weights[1235] <= 185;
		weights[1236] <= 59;
		weights[1237] <= 89;
		weights[1238] <= 196;
		weights[1239] <= 197;
		weights[1240] <= 152;
		weights[1241] <= 139;
		weights[1242] <= 47;
		weights[1243] <= 245;
		weights[1244] <= 204;
		weights[1245] <= 150;
		weights[1246] <= 27;
		weights[1247] <= 201;
		weights[1248] <= 67;
		weights[1249] <= 176;
		weights[1250] <= 119;
		weights[1251] <= 139;
		weights[1252] <= 135;
		weights[1253] <= 38;
		weights[1254] <= 222;
		weights[1255] <= 32;
		weights[1256] <= 6;
		weights[1257] <= 12;
		weights[1258] <= 133;
		weights[1259] <= 180;
		weights[1260] <= 48;
		weights[1261] <= 134;
		weights[1262] <= 255;
		weights[1263] <= 242;
		weights[1264] <= 11;
		weights[1265] <= 129;
		weights[1266] <= 133;
		weights[1267] <= 139;
		weights[1268] <= 158;
		weights[1269] <= 254;
		weights[1270] <= 94;
		weights[1271] <= 81;
		weights[1272] <= 31;
		weights[1273] <= 106;
		weights[1274] <= 116;
		weights[1275] <= 119;
		weights[1276] <= 10;
		weights[1277] <= 93;
		weights[1278] <= 93;
		weights[1279] <= 219;
		weights[1280] <= 78;
		weights[1281] <= 102;
		weights[1282] <= 70;
		weights[1283] <= 194;
		weights[1284] <= 214;
		weights[1285] <= 185;
		weights[1286] <= 229;
		weights[1287] <= 212;
		weights[1288] <= 184;
		weights[1289] <= 44;
		weights[1290] <= 77;
		weights[1291] <= 119;
		weights[1292] <= 64;
		weights[1293] <= 122;
		weights[1294] <= 185;
		weights[1295] <= 222;
		weights[1296] <= 187;
		weights[1297] <= 154;
		weights[1298] <= 14;
		weights[1299] <= 13;
		weights[1300] <= 53;
		weights[1301] <= 78;
		weights[1302] <= 84;
		weights[1303] <= 99;
		weights[1304] <= 27;
		weights[1305] <= 161;
		weights[1306] <= 17;
		weights[1307] <= 82;
		weights[1308] <= 178;
		weights[1309] <= 80;
		weights[1310] <= 233;
		weights[1311] <= 235;
		weights[1312] <= 234;
		weights[1313] <= 157;
		weights[1314] <= 125;
		weights[1315] <= 62;
		weights[1316] <= 185;
		weights[1317] <= 184;
		weights[1318] <= 145;
		weights[1319] <= 108;
		weights[1320] <= 96;
		weights[1321] <= 229;
		weights[1322] <= 196;
		weights[1323] <= 45;
		weights[1324] <= 65;
		weights[1325] <= 198;
		weights[1326] <= 70;
		weights[1327] <= 134;
		weights[1328] <= 148;
		weights[1329] <= 53;
		weights[1330] <= 254;
		weights[1331] <= 29;
		weights[1332] <= 203;
		weights[1333] <= 88;
		weights[1334] <= 7;
		weights[1335] <= 128;
		weights[1336] <= 247;
		weights[1337] <= 84;
		weights[1338] <= 216;
		weights[1339] <= 239;
		weights[1340] <= 151;
		weights[1341] <= 236;
		weights[1342] <= 249;
		weights[1343] <= 128;
		weights[1344] <= 235;
		weights[1345] <= 11;
		weights[1346] <= 29;
		weights[1347] <= 183;
		weights[1348] <= 228;
		weights[1349] <= 97;
		weights[1350] <= 52;
		weights[1351] <= 235;
		weights[1352] <= 48;
		weights[1353] <= 242;
		weights[1354] <= 158;
		weights[1355] <= 136;
		weights[1356] <= 117;
		weights[1357] <= 211;
		weights[1358] <= 22;
		weights[1359] <= 210;
		weights[1360] <= 226;
		weights[1361] <= 222;
		weights[1362] <= 121;
		weights[1363] <= 49;
		weights[1364] <= 128;
		weights[1365] <= 194;
		weights[1366] <= 95;
		weights[1367] <= 13;
		weights[1368] <= 233;
		weights[1369] <= 92;
		weights[1370] <= 100;
		weights[1371] <= 120;
		weights[1372] <= 134;
		weights[1373] <= 138;
		weights[1374] <= 188;
		weights[1375] <= 26;
		weights[1376] <= 108;
		weights[1377] <= 159;
		weights[1378] <= 130;
		weights[1379] <= 179;
		weights[1380] <= 139;
		weights[1381] <= 183;
		weights[1382] <= 65;
		weights[1383] <= 112;
		weights[1384] <= 4;
		weights[1385] <= 140;
		weights[1386] <= 200;
		weights[1387] <= 32;
		weights[1388] <= 102;
		weights[1389] <= 61;
		weights[1390] <= 188;
		weights[1391] <= 85;
		weights[1392] <= 211;
		weights[1393] <= 20;
		weights[1394] <= 29;
		weights[1395] <= 134;
		weights[1396] <= 154;
		weights[1397] <= 169;
		weights[1398] <= 3;
		weights[1399] <= 81;
		weights[1400] <= 10;
		weights[1401] <= 247;
		weights[1402] <= 147;
		weights[1403] <= 9;
		weights[1404] <= 60;
		weights[1405] <= 26;
		weights[1406] <= 153;
		weights[1407] <= 167;
		weights[1408] <= 220;
		weights[1409] <= 136;
		weights[1410] <= 124;
		weights[1411] <= 77;
		weights[1412] <= 237;
		weights[1413] <= 198;
		weights[1414] <= 184;
		weights[1415] <= 124;
		weights[1416] <= 208;
		weights[1417] <= 250;
		weights[1418] <= 130;
		weights[1419] <= 127;
		weights[1420] <= 83;
		weights[1421] <= 62;
		weights[1422] <= 69;
		weights[1423] <= 52;
		weights[1424] <= 199;
		weights[1425] <= 195;
		weights[1426] <= 74;
		weights[1427] <= 60;
		weights[1428] <= 66;
		weights[1429] <= 80;
		weights[1430] <= 179;
		weights[1431] <= 37;
		weights[1432] <= 162;
		weights[1433] <= 224;
		weights[1434] <= 224;
		weights[1435] <= 132;
		weights[1436] <= 233;
		weights[1437] <= 231;
		weights[1438] <= 186;
		weights[1439] <= 237;
		weights[1440] <= 96;
		weights[1441] <= 241;
		weights[1442] <= 132;
		weights[1443] <= 56;
		weights[1444] <= 175;
		weights[1445] <= 206;
		weights[1446] <= 20;
		weights[1447] <= 166;
		weights[1448] <= 94;
		weights[1449] <= 174;
		weights[1450] <= 52;
		weights[1451] <= 154;
		weights[1452] <= 150;
		weights[1453] <= 185;
		weights[1454] <= 58;
		weights[1455] <= 219;
		weights[1456] <= 178;
		weights[1457] <= 205;
		weights[1458] <= 93;
		weights[1459] <= 143;
		weights[1460] <= 165;
		weights[1461] <= 148;
		weights[1462] <= 53;
		weights[1463] <= 191;
		weights[1464] <= 3;
		weights[1465] <= 103;
		weights[1466] <= 221;
		weights[1467] <= 4;
		weights[1468] <= 123;
		weights[1469] <= 15;
		weights[1470] <= 76;
		weights[1471] <= 150;
		weights[1472] <= 94;
		weights[1473] <= 3;
		weights[1474] <= 47;
		weights[1475] <= 65;
		weights[1476] <= 242;
		weights[1477] <= 120;
		weights[1478] <= 79;
		weights[1479] <= 25;
		weights[1480] <= 70;
		weights[1481] <= 17;
		weights[1482] <= 142;
		weights[1483] <= 12;
		weights[1484] <= 181;
		weights[1485] <= 96;
		weights[1486] <= 101;
		weights[1487] <= 83;
		weights[1488] <= 215;
		weights[1489] <= 236;
		weights[1490] <= 110;
		weights[1491] <= 145;
		weights[1492] <= 10;
		weights[1493] <= 206;
		weights[1494] <= 255;
		weights[1495] <= 242;
		weights[1496] <= 109;
		weights[1497] <= 18;
		weights[1498] <= 209;
		weights[1499] <= 29;
		weights[1500] <= 214;
		weights[1501] <= 29;
		weights[1502] <= 71;
		weights[1503] <= 48;
		weights[1504] <= 106;
		weights[1505] <= 255;
		weights[1506] <= 176;
		weights[1507] <= 52;
		weights[1508] <= 30;
		weights[1509] <= 175;
		weights[1510] <= 58;
		weights[1511] <= 64;
		weights[1512] <= 192;
		weights[1513] <= 193;
		weights[1514] <= 89;
		weights[1515] <= 140;
		weights[1516] <= 76;
		weights[1517] <= 64;
		weights[1518] <= 126;
		weights[1519] <= 32;
		weights[1520] <= 155;
		weights[1521] <= 119;
		weights[1522] <= 6;
		weights[1523] <= 201;
		weights[1524] <= 162;
		weights[1525] <= 227;
		weights[1526] <= 210;
		weights[1527] <= 59;
		weights[1528] <= 96;
		weights[1529] <= 232;
		weights[1530] <= 248;
		weights[1531] <= 217;
		weights[1532] <= 122;
		weights[1533] <= 149;
		weights[1534] <= 253;
		weights[1535] <= 50;
		weights[1536] <= 227;
		weights[1537] <= 121;
		weights[1538] <= 255;
		weights[1539] <= 39;
		weights[1540] <= 122;
		weights[1541] <= 20;
		weights[1542] <= 129;
		weights[1543] <= 179;
		weights[1544] <= 116;
		weights[1545] <= 251;
		weights[1546] <= 203;
		weights[1547] <= 67;
		weights[1548] <= 90;
		weights[1549] <= 121;
		weights[1550] <= 220;
		weights[1551] <= 183;
		weights[1552] <= 179;
		weights[1553] <= 67;
		weights[1554] <= 218;
		weights[1555] <= 94;
		weights[1556] <= 16;
		weights[1557] <= 88;
		weights[1558] <= 110;
		weights[1559] <= 211;
		weights[1560] <= 127;
		weights[1561] <= 30;
		weights[1562] <= 40;
		weights[1563] <= 185;
		weights[1564] <= 142;
		weights[1565] <= 87;
		weights[1566] <= 221;
		weights[1567] <= 120;
		weights[1568] <= 151;
		weights[1569] <= 81;
		weights[1570] <= 76;
		weights[1571] <= 146;
		weights[1572] <= 56;
		weights[1573] <= 166;
		weights[1574] <= 114;
		weights[1575] <= 94;
		weights[1576] <= 132;
		weights[1577] <= 199;
		weights[1578] <= 217;
		weights[1579] <= 206;
		weights[1580] <= 27;
		weights[1581] <= 250;
		weights[1582] <= 71;
		weights[1583] <= 193;
		weights[1584] <= 12;
		weights[1585] <= 155;
		weights[1586] <= 243;
		weights[1587] <= 10;
		weights[1588] <= 212;
		weights[1589] <= 203;
		weights[1590] <= 12;
		weights[1591] <= 41;
		weights[1592] <= 214;
		weights[1593] <= 190;
		weights[1594] <= 113;
		weights[1595] <= 18;
		weights[1596] <= 124;
		weights[1597] <= 187;
		weights[1598] <= 86;
		weights[1599] <= 158;
		weights[1600] <= 30;
		weights[1601] <= 158;
		weights[1602] <= 103;
		weights[1603] <= 29;
		weights[1604] <= 112;
		weights[1605] <= 64;
		weights[1606] <= 96;
		weights[1607] <= 110;
		weights[1608] <= 232;
		weights[1609] <= 236;
		weights[1610] <= 190;
		weights[1611] <= 153;
		weights[1612] <= 172;
		weights[1613] <= 106;
		weights[1614] <= 184;
		weights[1615] <= 11;
		weights[1616] <= 248;
		weights[1617] <= 154;
		weights[1618] <= 209;
		weights[1619] <= 39;
		weights[1620] <= 154;
		weights[1621] <= 183;
		weights[1622] <= 131;
		weights[1623] <= 162;
		weights[1624] <= 172;
		weights[1625] <= 175;
		weights[1626] <= 140;
		weights[1627] <= 184;
		weights[1628] <= 19;
		weights[1629] <= 196;
		weights[1630] <= 110;
		weights[1631] <= 219;
		weights[1632] <= 138;
		weights[1633] <= 7;
		weights[1634] <= 119;
		weights[1635] <= 16;
		weights[1636] <= 8;
		weights[1637] <= 200;
		weights[1638] <= 77;
		weights[1639] <= 178;
		weights[1640] <= 188;
		weights[1641] <= 153;
		weights[1642] <= 63;
		weights[1643] <= 175;
		weights[1644] <= 41;
		weights[1645] <= 130;
		weights[1646] <= 161;
		weights[1647] <= 178;
		weights[1648] <= 233;
		weights[1649] <= 120;
		weights[1650] <= 134;
		weights[1651] <= 88;
		weights[1652] <= 164;
		weights[1653] <= 94;
		weights[1654] <= 81;
		weights[1655] <= 124;
		weights[1656] <= 45;
		weights[1657] <= 156;
		weights[1658] <= 61;
		weights[1659] <= 232;
		weights[1660] <= 239;
		weights[1661] <= 33;
		weights[1662] <= 194;
		weights[1663] <= 192;
		weights[1664] <= 150;
		weights[1665] <= 140;
		weights[1666] <= 246;
		weights[1667] <= 244;
		weights[1668] <= 22;
		weights[1669] <= 227;
		weights[1670] <= 221;
		weights[1671] <= 210;
		weights[1672] <= 144;
		weights[1673] <= 253;
		weights[1674] <= 70;
		weights[1675] <= 129;
		weights[1676] <= 143;
		weights[1677] <= 51;
		weights[1678] <= 115;
		weights[1679] <= 203;
		weights[1680] <= 143;
		weights[1681] <= 248;
		weights[1682] <= 13;
		weights[1683] <= 122;
		weights[1684] <= 235;
		weights[1685] <= 253;
		weights[1686] <= 166;
		weights[1687] <= 213;
		weights[1688] <= 118;
		weights[1689] <= 184;
		weights[1690] <= 103;
		weights[1691] <= 136;
		weights[1692] <= 204;
		weights[1693] <= 250;
		weights[1694] <= 137;
		weights[1695] <= 171;
		weights[1696] <= 238;
		weights[1697] <= 92;
		weights[1698] <= 185;
		weights[1699] <= 203;
		weights[1700] <= 8;
		weights[1701] <= 72;
		weights[1702] <= 175;
		weights[1703] <= 135;
		weights[1704] <= 150;
		weights[1705] <= 140;
		weights[1706] <= 84;
		weights[1707] <= 6;
		weights[1708] <= 197;
		weights[1709] <= 252;
		weights[1710] <= 252;
		weights[1711] <= 118;
		weights[1712] <= 144;
		weights[1713] <= 156;
		weights[1714] <= 158;
		weights[1715] <= 211;
		weights[1716] <= 141;
		weights[1717] <= 208;
		weights[1718] <= 201;
		weights[1719] <= 156;
		weights[1720] <= 98;
		weights[1721] <= 109;
		weights[1722] <= 176;
		weights[1723] <= 72;
		weights[1724] <= 161;
		weights[1725] <= 218;
		weights[1726] <= 68;
		weights[1727] <= 218;
		weights[1728] <= 130;
		weights[1729] <= 143;
		weights[1730] <= 242;
		weights[1731] <= 150;
		weights[1732] <= 56;
		weights[1733] <= 154;
		weights[1734] <= 184;
		weights[1735] <= 163;
		weights[1736] <= 196;
		weights[1737] <= 27;
		weights[1738] <= 235;
		weights[1739] <= 50;
		weights[1740] <= 138;
		weights[1741] <= 12;
		weights[1742] <= 110;
		weights[1743] <= 227;
		weights[1744] <= 66;
		weights[1745] <= 104;
		weights[1746] <= 67;
		weights[1747] <= 179;
		weights[1748] <= 178;
		weights[1749] <= 251;
		weights[1750] <= 227;
		weights[1751] <= 91;
		weights[1752] <= 163;
		weights[1753] <= 195;
		weights[1754] <= 68;
		weights[1755] <= 230;
		weights[1756] <= 53;
		weights[1757] <= 99;
		weights[1758] <= 66;
		weights[1759] <= 68;
		weights[1760] <= 143;
		weights[1761] <= 119;
		weights[1762] <= 37;
		weights[1763] <= 41;
		weights[1764] <= 59;
		weights[1765] <= 33;
		weights[1766] <= 212;
		weights[1767] <= 10;
		weights[1768] <= 247;
		weights[1769] <= 147;
		weights[1770] <= 218;
		weights[1771] <= 48;
		weights[1772] <= 195;
		weights[1773] <= 253;
		weights[1774] <= 129;
		weights[1775] <= 251;
		weights[1776] <= 255;
		weights[1777] <= 82;
		weights[1778] <= 223;
		weights[1779] <= 75;
		weights[1780] <= 134;
		weights[1781] <= 207;
		weights[1782] <= 113;
		weights[1783] <= 151;
		weights[1784] <= 51;
		weights[1785] <= 37;
		weights[1786] <= 192;
		weights[1787] <= 212;
		weights[1788] <= 81;
		weights[1789] <= 66;
		weights[1790] <= 211;
		weights[1791] <= 159;
		weights[1792] <= 27;
		weights[1793] <= 28;
		weights[1794] <= 246;
		weights[1795] <= 182;
		weights[1796] <= 195;
		weights[1797] <= 93;
		weights[1798] <= 230;
		weights[1799] <= 134;
		weights[1800] <= 78;
		weights[1801] <= 178;
		weights[1802] <= 198;
		weights[1803] <= 71;
		weights[1804] <= 166;
		weights[1805] <= 242;
		weights[1806] <= 4;
		weights[1807] <= 246;
		weights[1808] <= 215;
		weights[1809] <= 100;
		weights[1810] <= 215;
		weights[1811] <= 83;
		weights[1812] <= 175;
		weights[1813] <= 184;
		weights[1814] <= 204;
		weights[1815] <= 103;
		weights[1816] <= 156;
		weights[1817] <= 138;
		weights[1818] <= 153;
		weights[1819] <= 139;
		weights[1820] <= 190;
		weights[1821] <= 139;
		weights[1822] <= 37;
		weights[1823] <= 219;
		weights[1824] <= 245;
		weights[1825] <= 238;
		weights[1826] <= 247;
		weights[1827] <= 128;
		weights[1828] <= 146;
		weights[1829] <= 207;
		weights[1830] <= 60;
		weights[1831] <= 150;
		weights[1832] <= 75;
		weights[1833] <= 121;
		weights[1834] <= 245;
		weights[1835] <= 155;
		weights[1836] <= 150;
		weights[1837] <= 242;
		weights[1838] <= 228;
		weights[1839] <= 132;
		weights[1840] <= 27;
		weights[1841] <= 205;
		weights[1842] <= 21;
		weights[1843] <= 202;
		weights[1844] <= 26;
		weights[1845] <= 179;
		weights[1846] <= 6;
		weights[1847] <= 142;
		weights[1848] <= 120;
		weights[1849] <= 29;
		weights[1850] <= 197;
		weights[1851] <= 245;
		weights[1852] <= 196;
		weights[1853] <= 116;
		weights[1854] <= 91;
		weights[1855] <= 70;
		weights[1856] <= 9;
		weights[1857] <= 141;
		weights[1858] <= 113;
		weights[1859] <= 70;
		weights[1860] <= 131;
		weights[1861] <= 74;
		weights[1862] <= 180;
		weights[1863] <= 71;
		weights[1864] <= 143;
		weights[1865] <= 157;
		weights[1866] <= 75;
		weights[1867] <= 10;
		weights[1868] <= 152;
		weights[1869] <= 91;
		weights[1870] <= 45;
		weights[1871] <= 212;
		weights[1872] <= 236;
		weights[1873] <= 20;
		weights[1874] <= 32;
		weights[1875] <= 246;
		weights[1876] <= 83;
		weights[1877] <= 83;
		weights[1878] <= 68;
		weights[1879] <= 91;
		weights[1880] <= 130;
		weights[1881] <= 32;
		weights[1882] <= 107;
		weights[1883] <= 58;
		weights[1884] <= 107;
		weights[1885] <= 66;
		weights[1886] <= 105;
		weights[1887] <= 90;
		weights[1888] <= 230;
		weights[1889] <= 45;
		weights[1890] <= 151;
		weights[1891] <= 21;
		weights[1892] <= 144;
		weights[1893] <= 33;
		weights[1894] <= 197;
		weights[1895] <= 27;
		weights[1896] <= 132;
		weights[1897] <= 72;
		weights[1898] <= 212;
		weights[1899] <= 219;
		weights[1900] <= 240;
		weights[1901] <= 68;
		weights[1902] <= 194;
		weights[1903] <= 42;
		weights[1904] <= 35;
		weights[1905] <= 197;
		weights[1906] <= 133;
		weights[1907] <= 38;
		weights[1908] <= 99;
		weights[1909] <= 238;
		weights[1910] <= 69;
		weights[1911] <= 57;
		weights[1912] <= 6;
		weights[1913] <= 254;
		weights[1914] <= 140;
		weights[1915] <= 141;
		weights[1916] <= 112;
		weights[1917] <= 201;
		weights[1918] <= 182;
		weights[1919] <= 184;
		weights[1920] <= 97;
		weights[1921] <= 46;
		weights[1922] <= 205;
		weights[1923] <= 202;
		weights[1924] <= 74;
		weights[1925] <= 250;
		weights[1926] <= 206;
		weights[1927] <= 133;
		weights[1928] <= 235;
		weights[1929] <= 93;
		weights[1930] <= 89;
		weights[1931] <= 93;
		weights[1932] <= 6;
		weights[1933] <= 79;
		weights[1934] <= 65;
		weights[1935] <= 204;
		weights[1936] <= 248;
		weights[1937] <= 161;
		weights[1938] <= 211;
		weights[1939] <= 17;
		weights[1940] <= 241;
		weights[1941] <= 31;
		weights[1942] <= 32;
		weights[1943] <= 172;
		weights[1944] <= 34;
		weights[1945] <= 104;
		weights[1946] <= 145;
		weights[1947] <= 228;
		weights[1948] <= 130;
		weights[1949] <= 150;
		weights[1950] <= 85;
		weights[1951] <= 139;
		weights[1952] <= 90;
		weights[1953] <= 163;
		weights[1954] <= 126;
		weights[1955] <= 129;
		weights[1956] <= 16;
		weights[1957] <= 146;
		weights[1958] <= 28;
		weights[1959] <= 2;
		weights[1960] <= 19;
		weights[1961] <= 8;
		weights[1962] <= 49;
		weights[1963] <= 50;
		weights[1964] <= 171;
		weights[1965] <= 33;
		weights[1966] <= 1;
		weights[1967] <= 54;
		weights[1968] <= 4;
		weights[1969] <= 115;
		weights[1970] <= 60;
		weights[1971] <= 222;
		weights[1972] <= 107;
		weights[1973] <= 76;
		weights[1974] <= 4;
		weights[1975] <= 182;
		weights[1976] <= 182;
		weights[1977] <= 254;
		weights[1978] <= 110;
		weights[1979] <= 235;
		weights[1980] <= 14;
		weights[1981] <= 208;
		weights[1982] <= 52;
		weights[1983] <= 180;
		weights[1984] <= 169;
		weights[1985] <= 171;
		weights[1986] <= 192;
		weights[1987] <= 55;
		weights[1988] <= 240;
		weights[1989] <= 72;
		weights[1990] <= 242;
		weights[1991] <= 109;
		weights[1992] <= 144;
		weights[1993] <= 151;
		weights[1994] <= 17;
		weights[1995] <= 227;
		weights[1996] <= 252;
		weights[1997] <= 133;
		weights[1998] <= 31;
		weights[1999] <= 88;
		weights[2000] <= 49;
		weights[2001] <= 63;
		weights[2002] <= 107;
		weights[2003] <= 124;
		weights[2004] <= 102;
		weights[2005] <= 164;
		weights[2006] <= 12;
		weights[2007] <= 114;
		weights[2008] <= 80;
		weights[2009] <= 89;
		weights[2010] <= 164;
		weights[2011] <= 211;
		weights[2012] <= 65;
		weights[2013] <= 97;
		weights[2014] <= 250;
		weights[2015] <= 212;
		weights[2016] <= 19;
		weights[2017] <= 235;
		weights[2018] <= 69;
		weights[2019] <= 152;
		weights[2020] <= 21;
		weights[2021] <= 235;
		weights[2022] <= 232;
		weights[2023] <= 116;
		weights[2024] <= 155;
		weights[2025] <= 247;
		weights[2026] <= 247;
		weights[2027] <= 250;
		weights[2028] <= 216;
		weights[2029] <= 7;
		weights[2030] <= 15;
		weights[2031] <= 218;
		weights[2032] <= 125;
		weights[2033] <= 49;
		weights[2034] <= 139;
		weights[2035] <= 77;
		weights[2036] <= 61;
		weights[2037] <= 180;
		weights[2038] <= 249;
		weights[2039] <= 75;
		weights[2040] <= 240;
		weights[2041] <= 159;
		weights[2042] <= 238;
		weights[2043] <= 20;
		weights[2044] <= 87;
		weights[2045] <= 236;
		weights[2046] <= 44;
		weights[2047] <= 181;
		weights[2048] <= 209;
		weights[2049] <= 168;
		weights[2050] <= 8;
		weights[2051] <= 11;
		weights[2052] <= 149;
		weights[2053] <= 9;
		weights[2054] <= 146;
		weights[2055] <= 105;
		weights[2056] <= 52;
		weights[2057] <= 123;
		weights[2058] <= 66;
		weights[2059] <= 83;
		weights[2060] <= 203;
		weights[2061] <= 168;
		weights[2062] <= 32;
		weights[2063] <= 113;
		weights[2064] <= 195;
		weights[2065] <= 67;
		weights[2066] <= 101;
		weights[2067] <= 79;
		weights[2068] <= 92;
		weights[2069] <= 195;
		weights[2070] <= 53;
		weights[2071] <= 103;
		weights[2072] <= 13;
		weights[2073] <= 227;
		weights[2074] <= 8;
		weights[2075] <= 3;
		weights[2076] <= 219;
		weights[2077] <= 204;
		weights[2078] <= 177;
		weights[2079] <= 13;
		weights[2080] <= 50;
		weights[2081] <= 248;
		weights[2082] <= 18;
		weights[2083] <= 28;
		weights[2084] <= 52;
		weights[2085] <= 179;
		weights[2086] <= 50;
		weights[2087] <= 242;
		weights[2088] <= 8;
		weights[2089] <= 117;
		weights[2090] <= 32;
		weights[2091] <= 144;
		weights[2092] <= 3;
		weights[2093] <= 37;
		weights[2094] <= 110;
		weights[2095] <= 116;
		weights[2096] <= 87;
		weights[2097] <= 153;
		weights[2098] <= 4;
		weights[2099] <= 22;
		weights[2100] <= 91;
		weights[2101] <= 125;
		weights[2102] <= 178;
		weights[2103] <= 112;
		weights[2104] <= 164;
		weights[2105] <= 82;
		weights[2106] <= 156;
		weights[2107] <= 27;
		weights[2108] <= 199;
		weights[2109] <= 57;
		weights[2110] <= 69;
		weights[2111] <= 80;
		weights[2112] <= 131;
		weights[2113] <= 184;
		weights[2114] <= 147;
		weights[2115] <= 69;
		weights[2116] <= 119;
		weights[2117] <= 171;
		weights[2118] <= 46;
		weights[2119] <= 248;
		weights[2120] <= 235;
		weights[2121] <= 129;
		weights[2122] <= 69;
		weights[2123] <= 5;
		weights[2124] <= 71;
		weights[2125] <= 19;
		weights[2126] <= 133;
		weights[2127] <= 134;
		weights[2128] <= 3;
		weights[2129] <= 45;
		weights[2130] <= 220;
		weights[2131] <= 100;
		weights[2132] <= 7;
		weights[2133] <= 226;
		weights[2134] <= 155;
		weights[2135] <= 166;
		weights[2136] <= 243;
		weights[2137] <= 125;
		weights[2138] <= 104;
		weights[2139] <= 210;
		weights[2140] <= 131;
		weights[2141] <= 39;
		weights[2142] <= 155;
		weights[2143] <= 167;
		weights[2144] <= 50;
		weights[2145] <= 204;
		weights[2146] <= 166;
		weights[2147] <= 217;
		weights[2148] <= 166;
		weights[2149] <= 29;
		weights[2150] <= 138;
		weights[2151] <= 31;
		weights[2152] <= 111;
		weights[2153] <= 42;
		weights[2154] <= 98;
		weights[2155] <= 218;
		weights[2156] <= 192;
		weights[2157] <= 144;
		weights[2158] <= 39;
		weights[2159] <= 13;
		weights[2160] <= 69;
		weights[2161] <= 84;
		weights[2162] <= 92;
		weights[2163] <= 159;
		weights[2164] <= 238;
		weights[2165] <= 138;
		weights[2166] <= 216;
		weights[2167] <= 185;
		weights[2168] <= 34;
		weights[2169] <= 81;
		weights[2170] <= 5;
		weights[2171] <= 120;
		weights[2172] <= 156;
		weights[2173] <= 78;
		weights[2174] <= 74;
		weights[2175] <= 113;
		weights[2176] <= 250;
		weights[2177] <= 171;
		weights[2178] <= 55;
		weights[2179] <= 207;
		weights[2180] <= 43;
		weights[2181] <= 236;
		weights[2182] <= 211;
		weights[2183] <= 23;
		weights[2184] <= 150;
		weights[2185] <= 159;
		weights[2186] <= 126;
		weights[2187] <= 86;
		weights[2188] <= 179;
		weights[2189] <= 162;
		weights[2190] <= 195;
		weights[2191] <= 93;
		weights[2192] <= 134;
		weights[2193] <= 233;
		weights[2194] <= 202;
		weights[2195] <= 173;
		weights[2196] <= 218;
		weights[2197] <= 51;
		weights[2198] <= 201;
		weights[2199] <= 199;
		weights[2200] <= 111;
		weights[2201] <= 128;
		weights[2202] <= 47;
		weights[2203] <= 154;
		weights[2204] <= 50;
		weights[2205] <= 82;
		weights[2206] <= 85;
		weights[2207] <= 84;
		weights[2208] <= 1;
		weights[2209] <= 251;
		weights[2210] <= 78;
		weights[2211] <= 23;
		weights[2212] <= 151;
		weights[2213] <= 182;
		weights[2214] <= 28;
		weights[2215] <= 73;
		weights[2216] <= 213;
		weights[2217] <= 32;
		weights[2218] <= 217;
		weights[2219] <= 149;
		weights[2220] <= 35;
		weights[2221] <= 104;
		weights[2222] <= 210;
		weights[2223] <= 33;
		weights[2224] <= 36;
		weights[2225] <= 130;
		weights[2226] <= 193;
		weights[2227] <= 252;
		weights[2228] <= 99;
		weights[2229] <= 109;
		weights[2230] <= 132;
		weights[2231] <= 173;
		weights[2232] <= 110;
		weights[2233] <= 211;
		weights[2234] <= 136;
		weights[2235] <= 30;
		weights[2236] <= 163;
		weights[2237] <= 125;
		weights[2238] <= 45;
		weights[2239] <= 18;
		weights[2240] <= 7;
		weights[2241] <= 193;
		weights[2242] <= 10;
		weights[2243] <= 107;
		weights[2244] <= 19;
		weights[2245] <= 212;
		weights[2246] <= 32;
		weights[2247] <= 225;
		weights[2248] <= 153;
		weights[2249] <= 246;
		weights[2250] <= 60;
		weights[2251] <= 7;
		weights[2252] <= 80;
		weights[2253] <= 62;
		weights[2254] <= 61;
		weights[2255] <= 228;
		weights[2256] <= 120;
		weights[2257] <= 48;
		weights[2258] <= 186;
		weights[2259] <= 60;
		weights[2260] <= 219;
		weights[2261] <= 206;
		weights[2262] <= 246;
		weights[2263] <= 97;
		weights[2264] <= 126;
		weights[2265] <= 135;
		weights[2266] <= 114;
		weights[2267] <= 22;
		weights[2268] <= 217;
		weights[2269] <= 103;
		weights[2270] <= 16;
		weights[2271] <= 211;
		weights[2272] <= 148;
		weights[2273] <= 240;
		weights[2274] <= 239;
		weights[2275] <= 211;
		weights[2276] <= 197;
		weights[2277] <= 195;
		weights[2278] <= 95;
		weights[2279] <= 95;
		weights[2280] <= 230;
		weights[2281] <= 52;
		weights[2282] <= 240;
		weights[2283] <= 77;
		weights[2284] <= 249;
		weights[2285] <= 18;
		weights[2286] <= 147;
		weights[2287] <= 69;
		weights[2288] <= 137;
		weights[2289] <= 142;
		weights[2290] <= 251;
		weights[2291] <= 53;
		weights[2292] <= 246;
		weights[2293] <= 30;
		weights[2294] <= 222;
		weights[2295] <= 13;
		weights[2296] <= 101;
		weights[2297] <= 67;
		weights[2298] <= 204;
		weights[2299] <= 12;
		weights[2300] <= 4;
		weights[2301] <= 22;
		weights[2302] <= 3;
		weights[2303] <= 89;
		weights[2304] <= 138;
		weights[2305] <= 17;
		weights[2306] <= 7;
		weights[2307] <= 251;
		weights[2308] <= 237;
		weights[2309] <= 88;
		weights[2310] <= 254;
		weights[2311] <= 162;
		weights[2312] <= 132;
		weights[2313] <= 86;
		weights[2314] <= 213;
		weights[2315] <= 60;
		weights[2316] <= 85;
		weights[2317] <= 226;
		weights[2318] <= 20;
		weights[2319] <= 12;
		weights[2320] <= 158;
		weights[2321] <= 2;
		weights[2322] <= 120;
		weights[2323] <= 204;
		weights[2324] <= 43;
		weights[2325] <= 82;
		weights[2326] <= 21;
		weights[2327] <= 24;
		weights[2328] <= 231;
		weights[2329] <= 62;
		weights[2330] <= 230;
		weights[2331] <= 195;
		weights[2332] <= 124;
		weights[2333] <= 197;
		weights[2334] <= 172;
		weights[2335] <= 19;
		weights[2336] <= 216;
		weights[2337] <= 62;
		weights[2338] <= 111;
		weights[2339] <= 101;
		weights[2340] <= 77;
		weights[2341] <= 100;
		weights[2342] <= 56;
		weights[2343] <= 37;
		weights[2344] <= 74;
		weights[2345] <= 55;
		weights[2346] <= 195;
		weights[2347] <= 220;
		weights[2348] <= 83;
		weights[2349] <= 83;
		weights[2350] <= 252;
		weights[2351] <= 254;
		weights[2352] <= 72;
		weights[2353] <= 201;
		weights[2354] <= 53;
		weights[2355] <= 70;
		weights[2356] <= 88;
		weights[2357] <= 249;
		weights[2358] <= 18;
		weights[2359] <= 79;
		weights[2360] <= 184;
		weights[2361] <= 167;
		weights[2362] <= 150;
		weights[2363] <= 15;
		weights[2364] <= 161;
		weights[2365] <= 182;
		weights[2366] <= 143;
		weights[2367] <= 37;
		weights[2368] <= 221;
		weights[2369] <= 177;
		weights[2370] <= 24;
		weights[2371] <= 39;
		weights[2372] <= 164;
		weights[2373] <= 56;
		weights[2374] <= 241;
		weights[2375] <= 11;
		weights[2376] <= 113;
		weights[2377] <= 51;
		weights[2378] <= 212;
		weights[2379] <= 182;
		weights[2380] <= 41;
		weights[2381] <= 82;
		weights[2382] <= 114;
		weights[2383] <= 129;
		weights[2384] <= 59;
		weights[2385] <= 1;
		weights[2386] <= 245;
		weights[2387] <= 87;
		weights[2388] <= 179;
		weights[2389] <= 233;
		weights[2390] <= 126;
		weights[2391] <= 2;
		weights[2392] <= 112;
		weights[2393] <= 89;
		weights[2394] <= 82;
		weights[2395] <= 146;
		weights[2396] <= 134;
		weights[2397] <= 54;
		weights[2398] <= 208;
		weights[2399] <= 253;
		weights[2400] <= 232;
		weights[2401] <= 82;
		weights[2402] <= 141;
		weights[2403] <= 154;
		weights[2404] <= 219;
		weights[2405] <= 161;
		weights[2406] <= 101;
		weights[2407] <= 147;
		weights[2408] <= 180;
		weights[2409] <= 33;
		weights[2410] <= 103;
		weights[2411] <= 15;
		weights[2412] <= 202;
		weights[2413] <= 74;
		weights[2414] <= 99;
		weights[2415] <= 29;
		weights[2416] <= 171;
		weights[2417] <= 204;
		weights[2418] <= 102;
		weights[2419] <= 148;
		weights[2420] <= 51;
		weights[2421] <= 158;
		weights[2422] <= 21;
		weights[2423] <= 57;
		weights[2424] <= 146;
		weights[2425] <= 86;
		weights[2426] <= 20;
		weights[2427] <= 228;
		weights[2428] <= 33;
		weights[2429] <= 42;
		weights[2430] <= 159;
		weights[2431] <= 4;
		weights[2432] <= 153;
		weights[2433] <= 90;
		weights[2434] <= 97;
		weights[2435] <= 144;
		weights[2436] <= 97;
		weights[2437] <= 61;
		weights[2438] <= 146;
		weights[2439] <= 235;
		weights[2440] <= 135;
		weights[2441] <= 10;
		weights[2442] <= 235;
		weights[2443] <= 77;
		weights[2444] <= 205;
		weights[2445] <= 176;
		weights[2446] <= 219;
		weights[2447] <= 153;
		weights[2448] <= 149;
		weights[2449] <= 224;
		weights[2450] <= 205;
		weights[2451] <= 245;
		weights[2452] <= 239;
		weights[2453] <= 90;
		weights[2454] <= 48;
		weights[2455] <= 233;
		weights[2456] <= 232;
		weights[2457] <= 113;
		weights[2458] <= 10;
		weights[2459] <= 213;
		weights[2460] <= 233;
		weights[2461] <= 234;
		weights[2462] <= 12;
		weights[2463] <= 104;
		weights[2464] <= 81;
		weights[2465] <= 59;
		weights[2466] <= 51;
		weights[2467] <= 72;
		weights[2468] <= 216;
		weights[2469] <= 96;
		weights[2470] <= 227;
		weights[2471] <= 147;
		weights[2472] <= 178;
		weights[2473] <= 219;
		weights[2474] <= 2;
		weights[2475] <= 7;
		weights[2476] <= 61;
		weights[2477] <= 86;
		weights[2478] <= 68;
		weights[2479] <= 153;
		weights[2480] <= 195;
		weights[2481] <= 203;
		weights[2482] <= 128;
		weights[2483] <= 182;
		weights[2484] <= 86;
		weights[2485] <= 247;
		weights[2486] <= 225;
		weights[2487] <= 38;
		weights[2488] <= 95;
		weights[2489] <= 218;
		weights[2490] <= 158;
		weights[2491] <= 146;
		weights[2492] <= 19;
		weights[2493] <= 10;
		weights[2494] <= 89;
		weights[2495] <= 195;
		weights[2496] <= 53;
		weights[2497] <= 55;
		weights[2498] <= 110;
		weights[2499] <= 59;
		weights[2500] <= 174;
		weights[2501] <= 244;
		weights[2502] <= 154;
		weights[2503] <= 43;
		weights[2504] <= 15;
		weights[2505] <= 86;
		weights[2506] <= 131;
		weights[2507] <= 217;
		weights[2508] <= 89;
		weights[2509] <= 180;
		weights[2510] <= 207;
		weights[2511] <= 178;
		weights[2512] <= 163;
		weights[2513] <= 232;
		weights[2514] <= 91;
		weights[2515] <= 186;
		weights[2516] <= 117;
		weights[2517] <= 175;
		weights[2518] <= 195;
		weights[2519] <= 98;
		weights[2520] <= 74;
		weights[2521] <= 173;
		weights[2522] <= 253;
		weights[2523] <= 62;
		weights[2524] <= 201;
		weights[2525] <= 178;
		weights[2526] <= 60;
		weights[2527] <= 156;
		weights[2528] <= 145;
		weights[2529] <= 28;
		weights[2530] <= 94;
		weights[2531] <= 212;
		weights[2532] <= 20;
		weights[2533] <= 254;
		weights[2534] <= 224;
		weights[2535] <= 48;
		weights[2536] <= 13;
		weights[2537] <= 223;
		weights[2538] <= 17;
		weights[2539] <= 106;
		weights[2540] <= 152;
		weights[2541] <= 120;
		weights[2542] <= 60;
		weights[2543] <= 86;
		weights[2544] <= 242;
		weights[2545] <= 159;
		weights[2546] <= 137;
		weights[2547] <= 168;
		weights[2548] <= 47;
		weights[2549] <= 239;
		weights[2550] <= 2;
		weights[2551] <= 78;
		weights[2552] <= 25;
		weights[2553] <= 144;
		weights[2554] <= 146;
		weights[2555] <= 206;
		weights[2556] <= 118;
		weights[2557] <= 130;
		weights[2558] <= 230;
		weights[2559] <= 218;
		weights[2560] <= 60;
		weights[2561] <= 71;
		weights[2562] <= 68;
		weights[2563] <= 40;
		weights[2564] <= 41;
		weights[2565] <= 197;
		weights[2566] <= 115;
		weights[2567] <= 47;
		weights[2568] <= 112;
		weights[2569] <= 209;
		weights[2570] <= 215;
		weights[2571] <= 79;
		weights[2572] <= 199;
		weights[2573] <= 34;
		weights[2574] <= 65;
		weights[2575] <= 249;
		weights[2576] <= 243;
		weights[2577] <= 206;
		weights[2578] <= 61;
		weights[2579] <= 70;
		weights[2580] <= 232;
		weights[2581] <= 101;
		weights[2582] <= 152;
		weights[2583] <= 14;
		weights[2584] <= 40;
		weights[2585] <= 27;
		weights[2586] <= 113;
		weights[2587] <= 98;
		weights[2588] <= 136;
		weights[2589] <= 50;
		weights[2590] <= 134;
		weights[2591] <= 194;
		weights[2592] <= 154;
		weights[2593] <= 167;
		weights[2594] <= 50;
		weights[2595] <= 136;
		weights[2596] <= 13;
		weights[2597] <= 86;
		weights[2598] <= 49;
		weights[2599] <= 161;
		weights[2600] <= 144;
		weights[2601] <= 70;
		weights[2602] <= 133;
		weights[2603] <= 26;
		weights[2604] <= 116;
		weights[2605] <= 38;
		weights[2606] <= 173;
		weights[2607] <= 72;
		weights[2608] <= 199;
		weights[2609] <= 218;
		weights[2610] <= 234;
		weights[2611] <= 187;
		weights[2612] <= 77;
		weights[2613] <= 101;
		weights[2614] <= 69;
		weights[2615] <= 203;
		weights[2616] <= 186;
		weights[2617] <= 148;
		weights[2618] <= 124;
		weights[2619] <= 129;
		weights[2620] <= 219;
		weights[2621] <= 241;
		weights[2622] <= 213;
		weights[2623] <= 196;
		weights[2624] <= 246;
		weights[2625] <= 33;
		weights[2626] <= 22;
		weights[2627] <= 197;
		weights[2628] <= 50;
		weights[2629] <= 236;
		weights[2630] <= 157;
		weights[2631] <= 205;
		weights[2632] <= 178;
		weights[2633] <= 15;
		weights[2634] <= 230;
		weights[2635] <= 164;
		weights[2636] <= 241;
		weights[2637] <= 185;
		weights[2638] <= 146;
		weights[2639] <= 229;
		weights[2640] <= 24;
		weights[2641] <= 10;
		weights[2642] <= 140;
		weights[2643] <= 232;
		weights[2644] <= 140;
		weights[2645] <= 109;
		weights[2646] <= 253;
		weights[2647] <= 135;
		weights[2648] <= 198;
		weights[2649] <= 65;
		weights[2650] <= 30;
		weights[2651] <= 213;
		weights[2652] <= 150;
		weights[2653] <= 22;
		weights[2654] <= 136;
		weights[2655] <= 2;
		weights[2656] <= 78;
		weights[2657] <= 83;
		weights[2658] <= 227;
		weights[2659] <= 110;
		weights[2660] <= 39;
		weights[2661] <= 31;
		weights[2662] <= 196;
		weights[2663] <= 41;
		weights[2664] <= 77;
		weights[2665] <= 72;
		weights[2666] <= 187;
		weights[2667] <= 109;
		weights[2668] <= 58;
		weights[2669] <= 123;
		weights[2670] <= 224;
		weights[2671] <= 144;
		weights[2672] <= 50;
		weights[2673] <= 130;
		weights[2674] <= 230;
		weights[2675] <= 118;
		weights[2676] <= 11;
		weights[2677] <= 61;
		weights[2678] <= 59;
		weights[2679] <= 144;
		weights[2680] <= 5;
		weights[2681] <= 192;
		weights[2682] <= 83;
		weights[2683] <= 13;
		weights[2684] <= 192;
		weights[2685] <= 112;
		weights[2686] <= 231;
		weights[2687] <= 53;
		weights[2688] <= 90;
		weights[2689] <= 236;
		weights[2690] <= 32;
		weights[2691] <= 178;
		weights[2692] <= 180;
		weights[2693] <= 15;
		weights[2694] <= 183;
		weights[2695] <= 206;
		weights[2696] <= 155;
		weights[2697] <= 10;
		weights[2698] <= 75;
		weights[2699] <= 84;
		weights[2700] <= 97;
		weights[2701] <= 13;
		weights[2702] <= 62;
		weights[2703] <= 75;
		weights[2704] <= 50;
		weights[2705] <= 184;
		weights[2706] <= 152;
		weights[2707] <= 175;
		weights[2708] <= 78;
		weights[2709] <= 249;
		weights[2710] <= 67;
		weights[2711] <= 16;
		weights[2712] <= 198;
		weights[2713] <= 180;
		weights[2714] <= 61;
		weights[2715] <= 80;
		weights[2716] <= 218;
		weights[2717] <= 107;
		weights[2718] <= 174;
		weights[2719] <= 85;
		weights[2720] <= 140;
		weights[2721] <= 178;
		weights[2722] <= 26;
		weights[2723] <= 190;
		weights[2724] <= 80;
		weights[2725] <= 135;
		weights[2726] <= 69;
		weights[2727] <= 124;
		weights[2728] <= 65;
		weights[2729] <= 56;
		weights[2730] <= 162;
		weights[2731] <= 217;
		weights[2732] <= 194;
		weights[2733] <= 79;
		weights[2734] <= 180;
		weights[2735] <= 133;
		weights[2736] <= 239;
		weights[2737] <= 142;
		weights[2738] <= 94;
		weights[2739] <= 113;
		weights[2740] <= 50;
		weights[2741] <= 116;
		weights[2742] <= 200;
		weights[2743] <= 173;
		weights[2744] <= 107;
		weights[2745] <= 7;
		weights[2746] <= 36;
		weights[2747] <= 183;
		weights[2748] <= 46;
		weights[2749] <= 41;
		weights[2750] <= 211;
		weights[2751] <= 120;
		weights[2752] <= 154;
		weights[2753] <= 173;
		weights[2754] <= 92;
		weights[2755] <= 166;
		weights[2756] <= 58;
		weights[2757] <= 65;
		weights[2758] <= 94;
		weights[2759] <= 66;
		weights[2760] <= 96;
		weights[2761] <= 204;
		weights[2762] <= 107;
		weights[2763] <= 13;
		weights[2764] <= 161;
		weights[2765] <= 41;
		weights[2766] <= 96;
		weights[2767] <= 44;
		weights[2768] <= 105;
		weights[2769] <= 98;
		weights[2770] <= 228;
		weights[2771] <= 209;
		weights[2772] <= 236;
		weights[2773] <= 87;
		weights[2774] <= 153;
		weights[2775] <= 129;
		weights[2776] <= 61;
		weights[2777] <= 189;
		weights[2778] <= 119;
		weights[2779] <= 235;
		weights[2780] <= 35;
		weights[2781] <= 125;
		weights[2782] <= 65;
		weights[2783] <= 235;
		weights[2784] <= 79;
		weights[2785] <= 146;
		weights[2786] <= 70;
		weights[2787] <= 37;
		weights[2788] <= 159;
		weights[2789] <= 54;
		weights[2790] <= 24;
		weights[2791] <= 143;
		weights[2792] <= 21;
		weights[2793] <= 198;
		weights[2794] <= 58;
		weights[2795] <= 30;
		weights[2796] <= 11;
		weights[2797] <= 132;
		weights[2798] <= 140;
		weights[2799] <= 40;
		weights[2800] <= 216;
		weights[2801] <= 83;
		weights[2802] <= 61;
		weights[2803] <= 164;
		weights[2804] <= 57;
		weights[2805] <= 216;
		weights[2806] <= 27;
		weights[2807] <= 241;
		weights[2808] <= 9;
		weights[2809] <= 198;
		weights[2810] <= 191;
		weights[2811] <= 74;
		weights[2812] <= 184;
		weights[2813] <= 73;
		weights[2814] <= 195;
		weights[2815] <= 241;
		weights[2816] <= 1;
		weights[2817] <= 45;
		weights[2818] <= 70;
		weights[2819] <= 119;
		weights[2820] <= 41;
		weights[2821] <= 157;
		weights[2822] <= 64;
		weights[2823] <= 67;
		weights[2824] <= 103;
		weights[2825] <= 113;
		weights[2826] <= 31;
		weights[2827] <= 91;
		weights[2828] <= 48;
		weights[2829] <= 104;
		weights[2830] <= 20;
		weights[2831] <= 125;
		weights[2832] <= 166;
		weights[2833] <= 139;
		weights[2834] <= 38;
		weights[2835] <= 88;
		weights[2836] <= 51;
		weights[2837] <= 102;
		weights[2838] <= 127;
		weights[2839] <= 118;
		weights[2840] <= 177;
		weights[2841] <= 210;
		weights[2842] <= 234;
		weights[2843] <= 201;
		weights[2844] <= 76;
		weights[2845] <= 38;
		weights[2846] <= 68;
		weights[2847] <= 145;
		weights[2848] <= 37;
		weights[2849] <= 215;
		weights[2850] <= 197;
		weights[2851] <= 115;
		weights[2852] <= 36;
		weights[2853] <= 88;
		weights[2854] <= 42;
		weights[2855] <= 97;
		weights[2856] <= 114;
		weights[2857] <= 113;
		weights[2858] <= 208;
		weights[2859] <= 224;
		weights[2860] <= 180;
		weights[2861] <= 250;
		weights[2862] <= 36;
		weights[2863] <= 87;
		weights[2864] <= 242;
		weights[2865] <= 74;
		weights[2866] <= 39;
		weights[2867] <= 111;
		weights[2868] <= 157;
		weights[2869] <= 245;
		weights[2870] <= 170;
		weights[2871] <= 222;
		weights[2872] <= 170;
		weights[2873] <= 235;
		weights[2874] <= 143;
		weights[2875] <= 181;
		weights[2876] <= 12;
		weights[2877] <= 123;
		weights[2878] <= 108;
		weights[2879] <= 32;
		weights[2880] <= 153;
		weights[2881] <= 247;
		weights[2882] <= 250;
		weights[2883] <= 17;
		weights[2884] <= 89;
		weights[2885] <= 187;
		weights[2886] <= 121;
		weights[2887] <= 80;
		weights[2888] <= 243;
		weights[2889] <= 112;
		weights[2890] <= 50;
		weights[2891] <= 230;
		weights[2892] <= 39;
		weights[2893] <= 72;
		weights[2894] <= 103;
		weights[2895] <= 108;
		weights[2896] <= 89;
		weights[2897] <= 108;
		weights[2898] <= 163;
		weights[2899] <= 203;
		weights[2900] <= 25;
		weights[2901] <= 110;
		weights[2902] <= 164;
		weights[2903] <= 249;
		weights[2904] <= 112;
		weights[2905] <= 165;
		weights[2906] <= 156;
		weights[2907] <= 164;
		weights[2908] <= 215;
		weights[2909] <= 179;
		weights[2910] <= 7;
		weights[2911] <= 95;
		weights[2912] <= 51;
		weights[2913] <= 178;
		weights[2914] <= 204;
		weights[2915] <= 76;
		weights[2916] <= 69;
		weights[2917] <= 150;
		weights[2918] <= 232;
		weights[2919] <= 70;
		weights[2920] <= 59;
		weights[2921] <= 137;
		weights[2922] <= 8;
		weights[2923] <= 140;
		weights[2924] <= 160;
		weights[2925] <= 124;
		weights[2926] <= 84;
		weights[2927] <= 203;
		weights[2928] <= 84;
		weights[2929] <= 142;
		weights[2930] <= 26;
		weights[2931] <= 144;
		weights[2932] <= 160;
		weights[2933] <= 2;
		weights[2934] <= 2;
		weights[2935] <= 78;
		weights[2936] <= 101;
		weights[2937] <= 42;
		weights[2938] <= 104;
		weights[2939] <= 59;
		weights[2940] <= 33;
		weights[2941] <= 201;
		weights[2942] <= 150;
		weights[2943] <= 97;
		weights[2944] <= 106;
		weights[2945] <= 239;
		weights[2946] <= 38;
		weights[2947] <= 230;
		weights[2948] <= 227;
		weights[2949] <= 194;
		weights[2950] <= 224;
		weights[2951] <= 234;
		weights[2952] <= 156;
		weights[2953] <= 161;
		weights[2954] <= 58;
		weights[2955] <= 229;
		weights[2956] <= 154;
		weights[2957] <= 197;
		weights[2958] <= 25;
		weights[2959] <= 217;
		weights[2960] <= 94;
		weights[2961] <= 225;
		weights[2962] <= 142;
		weights[2963] <= 36;
		weights[2964] <= 59;
		weights[2965] <= 224;
		weights[2966] <= 126;
		weights[2967] <= 230;
		weights[2968] <= 140;
		weights[2969] <= 88;
		weights[2970] <= 115;
		weights[2971] <= 166;
		weights[2972] <= 63;
		weights[2973] <= 134;
		weights[2974] <= 129;
		weights[2975] <= 207;
		weights[2976] <= 37;
		weights[2977] <= 233;
		weights[2978] <= 251;
		weights[2979] <= 122;
		weights[2980] <= 66;
		weights[2981] <= 5;
		weights[2982] <= 230;
		weights[2983] <= 85;
		weights[2984] <= 251;
		weights[2985] <= 85;
		weights[2986] <= 50;
		weights[2987] <= 200;
		weights[2988] <= 60;
		weights[2989] <= 123;
		weights[2990] <= 171;
		weights[2991] <= 129;
		weights[2992] <= 202;
		weights[2993] <= 194;
		weights[2994] <= 158;
		weights[2995] <= 238;
		weights[2996] <= 168;
		weights[2997] <= 242;
		weights[2998] <= 137;
		weights[2999] <= 120;
		weights[3000] <= 234;
		weights[3001] <= 98;
		weights[3002] <= 14;
		weights[3003] <= 89;
		weights[3004] <= 68;
		weights[3005] <= 132;
		weights[3006] <= 8;
		weights[3007] <= 233;
		weights[3008] <= 26;
		weights[3009] <= 110;
		weights[3010] <= 36;
		weights[3011] <= 232;
		weights[3012] <= 234;
		weights[3013] <= 141;
		weights[3014] <= 239;
		weights[3015] <= 46;
		weights[3016] <= 6;
		weights[3017] <= 29;
		weights[3018] <= 55;
		weights[3019] <= 191;
		weights[3020] <= 135;
		weights[3021] <= 190;
		weights[3022] <= 12;
		weights[3023] <= 86;
		weights[3024] <= 107;
		weights[3025] <= 100;
		weights[3026] <= 216;
		weights[3027] <= 197;
		weights[3028] <= 119;
		weights[3029] <= 40;
		weights[3030] <= 136;
		weights[3031] <= 174;
		weights[3032] <= 65;
		weights[3033] <= 125;
		weights[3034] <= 167;
		weights[3035] <= 152;
		weights[3036] <= 81;
		weights[3037] <= 159;
		weights[3038] <= 244;
		weights[3039] <= 129;
		weights[3040] <= 183;
		weights[3041] <= 179;
		weights[3042] <= 216;
		weights[3043] <= 176;
		weights[3044] <= 136;
		weights[3045] <= 158;
		weights[3046] <= 5;
		weights[3047] <= 235;
		weights[3048] <= 63;
		weights[3049] <= 146;
		weights[3050] <= 5;
		weights[3051] <= 44;
		weights[3052] <= 136;
		weights[3053] <= 224;
		weights[3054] <= 104;
		weights[3055] <= 203;
		weights[3056] <= 59;
		weights[3057] <= 139;
		weights[3058] <= 32;
		weights[3059] <= 194;
		weights[3060] <= 168;
		weights[3061] <= 30;
		weights[3062] <= 113;
		weights[3063] <= 169;
		weights[3064] <= 72;
		weights[3065] <= 206;
		weights[3066] <= 38;
		weights[3067] <= 4;
		weights[3068] <= 195;
		weights[3069] <= 7;
		weights[3070] <= 95;
		weights[3071] <= 99;
		weights[3072] <= 9;
		weights[3073] <= 83;
		weights[3074] <= 99;
		weights[3075] <= 148;
		weights[3076] <= 212;
		weights[3077] <= 250;
		weights[3078] <= 1;
		weights[3079] <= 173;
		weights[3080] <= 205;
		weights[3081] <= 132;
		weights[3082] <= 98;
		weights[3083] <= 10;
		weights[3084] <= 69;
		weights[3085] <= 155;
		weights[3086] <= 14;
		weights[3087] <= 75;
		weights[3088] <= 251;
		weights[3089] <= 158;
		weights[3090] <= 117;
		weights[3091] <= 76;
		weights[3092] <= 8;
		weights[3093] <= 217;
		weights[3094] <= 167;
		weights[3095] <= 154;
		weights[3096] <= 3;
		weights[3097] <= 43;
		weights[3098] <= 190;
		weights[3099] <= 16;
		weights[3100] <= 77;
		weights[3101] <= 43;
		weights[3102] <= 27;
		weights[3103] <= 226;
		weights[3104] <= 103;
		weights[3105] <= 187;
		weights[3106] <= 79;
		weights[3107] <= 141;
		weights[3108] <= 37;
		weights[3109] <= 21;
		weights[3110] <= 171;
		weights[3111] <= 182;
		weights[3112] <= 226;
		weights[3113] <= 164;
		weights[3114] <= 67;
		weights[3115] <= 74;
		weights[3116] <= 47;
		weights[3117] <= 240;
		weights[3118] <= 113;
		weights[3119] <= 116;
		weights[3120] <= 165;
		weights[3121] <= 155;
		weights[3122] <= 133;
		weights[3123] <= 182;
		weights[3124] <= 102;
		weights[3125] <= 177;
		weights[3126] <= 29;
		weights[3127] <= 234;
		weights[3128] <= 215;
		weights[3129] <= 33;
		weights[3130] <= 42;
		weights[3131] <= 210;
		weights[3132] <= 221;
		weights[3133] <= 113;
		weights[3134] <= 206;
		weights[3135] <= 9;
		weights[3136] <= 156;
		weights[3137] <= 179;
		weights[3138] <= 28;
		weights[3139] <= 43;
		weights[3140] <= 118;
		weights[3141] <= 56;
		weights[3142] <= 167;
		weights[3143] <= 213;
		weights[3144] <= 42;
		weights[3145] <= 67;
		weights[3146] <= 30;
		weights[3147] <= 118;
		weights[3148] <= 78;
		weights[3149] <= 241;
		weights[3150] <= 86;
		weights[3151] <= 231;
		weights[3152] <= 174;
		weights[3153] <= 119;
		weights[3154] <= 240;
		weights[3155] <= 177;
		weights[3156] <= 191;
		weights[3157] <= 73;
		weights[3158] <= 73;
		weights[3159] <= 179;
		weights[3160] <= 3;
		weights[3161] <= 74;
		weights[3162] <= 176;
		weights[3163] <= 130;
		weights[3164] <= 19;
		weights[3165] <= 141;
		weights[3166] <= 110;
		weights[3167] <= 233;
		weights[3168] <= 247;
		weights[3169] <= 11;
		weights[3170] <= 63;
		weights[3171] <= 101;
		weights[3172] <= 212;
		weights[3173] <= 150;
		weights[3174] <= 28;
		weights[3175] <= 88;
		weights[3176] <= 84;
		weights[3177] <= 79;
		weights[3178] <= 73;
		weights[3179] <= 229;
		weights[3180] <= 210;
		weights[3181] <= 251;
		weights[3182] <= 24;
		weights[3183] <= 186;
		weights[3184] <= 92;
		weights[3185] <= 54;
		weights[3186] <= 96;
		weights[3187] <= 200;
		weights[3188] <= 208;
		weights[3189] <= 19;
		weights[3190] <= 140;
		weights[3191] <= 231;
		weights[3192] <= 81;
		weights[3193] <= 246;
		weights[3194] <= 125;
		weights[3195] <= 75;
		weights[3196] <= 20;
		weights[3197] <= 120;
		weights[3198] <= 190;
		weights[3199] <= 101;
		weights[3200] <= 205;
		weights[3201] <= 150;
		weights[3202] <= 170;
		weights[3203] <= 64;
		weights[3204] <= 223;
		weights[3205] <= 15;
		weights[3206] <= 120;
		weights[3207] <= 30;
		weights[3208] <= 227;
		weights[3209] <= 78;
		weights[3210] <= 2;
		weights[3211] <= 52;
		weights[3212] <= 201;
		weights[3213] <= 42;
		weights[3214] <= 126;
		weights[3215] <= 126;
		weights[3216] <= 38;
		weights[3217] <= 120;
		weights[3218] <= 82;
		weights[3219] <= 94;
		weights[3220] <= 239;
		weights[3221] <= 163;
		weights[3222] <= 227;
		weights[3223] <= 229;
		weights[3224] <= 94;
		weights[3225] <= 128;
		weights[3226] <= 189;
		weights[3227] <= 111;
		weights[3228] <= 21;
		weights[3229] <= 31;
		weights[3230] <= 133;
		weights[3231] <= 206;
		weights[3232] <= 119;
		weights[3233] <= 60;
		weights[3234] <= 236;
		weights[3235] <= 32;
		weights[3236] <= 27;
		weights[3237] <= 12;
		weights[3238] <= 154;
		weights[3239] <= 175;
		weights[3240] <= 135;
		weights[3241] <= 132;
		weights[3242] <= 147;
		weights[3243] <= 21;
		weights[3244] <= 71;
		weights[3245] <= 177;
		weights[3246] <= 46;
		weights[3247] <= 168;
		weights[3248] <= 92;
		weights[3249] <= 185;
		weights[3250] <= 125;
		weights[3251] <= 94;
		weights[3252] <= 123;
		weights[3253] <= 232;
		weights[3254] <= 171;
		weights[3255] <= 204;
		weights[3256] <= 53;
		weights[3257] <= 205;
		weights[3258] <= 230;
		weights[3259] <= 21;
		weights[3260] <= 238;
		weights[3261] <= 14;
		weights[3262] <= 79;
		weights[3263] <= 69;
		weights[3264] <= 105;
		weights[3265] <= 102;
		weights[3266] <= 102;
		weights[3267] <= 188;
		weights[3268] <= 116;
		weights[3269] <= 154;
		weights[3270] <= 74;
		weights[3271] <= 50;
		weights[3272] <= 13;
		weights[3273] <= 23;
		weights[3274] <= 114;
		weights[3275] <= 233;
		weights[3276] <= 148;
		weights[3277] <= 244;
		weights[3278] <= 228;
		weights[3279] <= 224;
		weights[3280] <= 203;
		weights[3281] <= 249;
		weights[3282] <= 124;
		weights[3283] <= 103;
		weights[3284] <= 86;
		weights[3285] <= 195;
		weights[3286] <= 91;
		weights[3287] <= 227;
		weights[3288] <= 17;
		weights[3289] <= 4;
		weights[3290] <= 66;
		weights[3291] <= 237;
		weights[3292] <= 69;
		weights[3293] <= 81;
		weights[3294] <= 65;
		weights[3295] <= 240;
		weights[3296] <= 144;
		weights[3297] <= 190;
		weights[3298] <= 139;
		weights[3299] <= 68;
		weights[3300] <= 110;
		weights[3301] <= 216;
		weights[3302] <= 46;
		weights[3303] <= 89;
		weights[3304] <= 8;
		weights[3305] <= 71;
		weights[3306] <= 152;
		weights[3307] <= 120;
		weights[3308] <= 210;
		weights[3309] <= 96;
		weights[3310] <= 247;
		weights[3311] <= 38;
		weights[3312] <= 83;
		weights[3313] <= 195;
		weights[3314] <= 127;
		weights[3315] <= 215;
		weights[3316] <= 249;
		weights[3317] <= 213;
		weights[3318] <= 119;
		weights[3319] <= 229;
		weights[3320] <= 41;
		weights[3321] <= 35;
		weights[3322] <= 29;
		weights[3323] <= 87;
		weights[3324] <= 168;
		weights[3325] <= 136;
		weights[3326] <= 255;
		weights[3327] <= 22;
		weights[3328] <= 63;
		weights[3329] <= 28;
		weights[3330] <= 166;
		weights[3331] <= 184;
		weights[3332] <= 241;
		weights[3333] <= 169;
		weights[3334] <= 152;
		weights[3335] <= 80;
		weights[3336] <= 136;
		weights[3337] <= 135;
		weights[3338] <= 7;
		weights[3339] <= 247;
		weights[3340] <= 224;
		weights[3341] <= 69;
		weights[3342] <= 25;
		weights[3343] <= 90;
		weights[3344] <= 128;
		weights[3345] <= 237;
		weights[3346] <= 37;
		weights[3347] <= 61;
		weights[3348] <= 22;
		weights[3349] <= 129;
		weights[3350] <= 135;
		weights[3351] <= 194;
		weights[3352] <= 81;
		weights[3353] <= 237;
		weights[3354] <= 172;
		weights[3355] <= 69;
		weights[3356] <= 52;
		weights[3357] <= 175;
		weights[3358] <= 31;
		weights[3359] <= 135;
		weights[3360] <= 70;
		weights[3361] <= 13;
		weights[3362] <= 178;
		weights[3363] <= 151;
		weights[3364] <= 208;
		weights[3365] <= 116;
		weights[3366] <= 119;
		weights[3367] <= 160;
		weights[3368] <= 85;
		weights[3369] <= 9;
		weights[3370] <= 97;
		weights[3371] <= 93;
		weights[3372] <= 199;
		weights[3373] <= 117;
		weights[3374] <= 154;
		weights[3375] <= 21;
		weights[3376] <= 249;
		weights[3377] <= 104;
		weights[3378] <= 237;
		weights[3379] <= 196;
		weights[3380] <= 213;
		weights[3381] <= 34;
		weights[3382] <= 205;
		weights[3383] <= 156;
		weights[3384] <= 163;
		weights[3385] <= 212;
		weights[3386] <= 81;
		weights[3387] <= 118;
		weights[3388] <= 37;
		weights[3389] <= 185;
		weights[3390] <= 182;
		weights[3391] <= 216;
		weights[3392] <= 206;
		weights[3393] <= 54;
		weights[3394] <= 227;
		weights[3395] <= 164;
		weights[3396] <= 254;
		weights[3397] <= 3;
		weights[3398] <= 188;
		weights[3399] <= 207;
		weights[3400] <= 164;
		weights[3401] <= 236;
		weights[3402] <= 22;
		weights[3403] <= 201;
		weights[3404] <= 212;
		weights[3405] <= 54;
		weights[3406] <= 106;
		weights[3407] <= 255;
		weights[3408] <= 13;
		weights[3409] <= 202;
		weights[3410] <= 4;
		weights[3411] <= 74;
		weights[3412] <= 58;
		weights[3413] <= 210;
		weights[3414] <= 35;
		weights[3415] <= 86;
		weights[3416] <= 236;
		weights[3417] <= 201;
		weights[3418] <= 52;
		weights[3419] <= 111;
		weights[3420] <= 123;
		weights[3421] <= 203;
		weights[3422] <= 211;
		weights[3423] <= 152;
		weights[3424] <= 250;
		weights[3425] <= 43;
		weights[3426] <= 206;
		weights[3427] <= 231;
		weights[3428] <= 27;
		weights[3429] <= 55;
		weights[3430] <= 251;
		weights[3431] <= 227;
		weights[3432] <= 137;
		weights[3433] <= 69;
		weights[3434] <= 213;
		weights[3435] <= 94;
		weights[3436] <= 246;
		weights[3437] <= 84;
		weights[3438] <= 1;
		weights[3439] <= 70;
		weights[3440] <= 166;
		weights[3441] <= 250;
		weights[3442] <= 115;
		weights[3443] <= 11;
		weights[3444] <= 245;
		weights[3445] <= 27;
		weights[3446] <= 239;
		weights[3447] <= 202;
		weights[3448] <= 47;
		weights[3449] <= 167;
		weights[3450] <= 11;
		weights[3451] <= 213;
		weights[3452] <= 239;
		weights[3453] <= 65;
		weights[3454] <= 195;
		weights[3455] <= 129;
		weights[3456] <= 207;
		weights[3457] <= 166;
		weights[3458] <= 14;
		weights[3459] <= 223;
		weights[3460] <= 185;
		weights[3461] <= 75;
		weights[3462] <= 134;
		weights[3463] <= 237;
		weights[3464] <= 225;
		weights[3465] <= 23;
		weights[3466] <= 128;
		weights[3467] <= 77;
		weights[3468] <= 130;
		weights[3469] <= 182;
		weights[3470] <= 168;
		weights[3471] <= 188;
		weights[3472] <= 241;
		weights[3473] <= 22;
		weights[3474] <= 35;
		weights[3475] <= 96;
		weights[3476] <= 240;
		weights[3477] <= 8;
		weights[3478] <= 197;
		weights[3479] <= 37;
		weights[3480] <= 145;
		weights[3481] <= 210;
		weights[3482] <= 175;
		weights[3483] <= 71;
		weights[3484] <= 180;
		weights[3485] <= 27;
		weights[3486] <= 17;
		weights[3487] <= 27;
		weights[3488] <= 5;
		weights[3489] <= 86;
		weights[3490] <= 125;
		weights[3491] <= 78;
		weights[3492] <= 21;
		weights[3493] <= 238;
		weights[3494] <= 92;
		weights[3495] <= 199;
		weights[3496] <= 65;
		weights[3497] <= 25;
		weights[3498] <= 18;
		weights[3499] <= 255;
		weights[3500] <= 155;
		weights[3501] <= 37;
		weights[3502] <= 219;
		weights[3503] <= 225;
		weights[3504] <= 16;
		weights[3505] <= 26;
		weights[3506] <= 193;
		weights[3507] <= 156;
		weights[3508] <= 128;
		weights[3509] <= 57;
		weights[3510] <= 175;
		weights[3511] <= 6;
		weights[3512] <= 235;
		weights[3513] <= 181;
		weights[3514] <= 28;
		weights[3515] <= 14;
		weights[3516] <= 219;
		weights[3517] <= 110;
		weights[3518] <= 101;
		weights[3519] <= 8;
		weights[3520] <= 11;
		weights[3521] <= 116;
		weights[3522] <= 95;
		weights[3523] <= 62;
		weights[3524] <= 228;
		weights[3525] <= 36;
		weights[3526] <= 92;
		weights[3527] <= 30;
		weights[3528] <= 98;
		weights[3529] <= 19;
		weights[3530] <= 135;
		weights[3531] <= 225;
		weights[3532] <= 182;
		weights[3533] <= 105;
		weights[3534] <= 254;
		weights[3535] <= 247;
		weights[3536] <= 22;
		weights[3537] <= 92;
		weights[3538] <= 121;
		weights[3539] <= 78;
		weights[3540] <= 191;
		weights[3541] <= 127;
		weights[3542] <= 113;
		weights[3543] <= 185;
		weights[3544] <= 68;
		weights[3545] <= 95;
		weights[3546] <= 190;
		weights[3547] <= 217;
		weights[3548] <= 91;
		weights[3549] <= 194;
		weights[3550] <= 33;
		weights[3551] <= 140;
		weights[3552] <= 158;
		weights[3553] <= 241;
		weights[3554] <= 79;
		weights[3555] <= 244;
		weights[3556] <= 192;
		weights[3557] <= 111;
		weights[3558] <= 203;
		weights[3559] <= 112;
		weights[3560] <= 234;
		weights[3561] <= 37;
		weights[3562] <= 25;
		weights[3563] <= 153;
		weights[3564] <= 149;
		weights[3565] <= 113;
		weights[3566] <= 153;
		weights[3567] <= 252;
		weights[3568] <= 245;
		weights[3569] <= 251;
		weights[3570] <= 44;
		weights[3571] <= 206;
		weights[3572] <= 81;
		weights[3573] <= 179;
		weights[3574] <= 145;
		weights[3575] <= 131;
		weights[3576] <= 78;
		weights[3577] <= 219;
		weights[3578] <= 95;
		weights[3579] <= 28;
		weights[3580] <= 205;
		weights[3581] <= 20;
		weights[3582] <= 30;
		weights[3583] <= 251;
		weights[3584] <= 13;
		weights[3585] <= 82;
		weights[3586] <= 154;
		weights[3587] <= 158;
		weights[3588] <= 98;
		weights[3589] <= 170;
		weights[3590] <= 208;
		weights[3591] <= 9;
		weights[3592] <= 247;
		weights[3593] <= 163;
		weights[3594] <= 29;
		weights[3595] <= 96;
		weights[3596] <= 252;
		weights[3597] <= 2;
		weights[3598] <= 96;
		weights[3599] <= 38;
		weights[3600] <= 175;
		weights[3601] <= 86;
		weights[3602] <= 220;
		weights[3603] <= 8;
		weights[3604] <= 20;
		weights[3605] <= 124;
		weights[3606] <= 55;
		weights[3607] <= 168;
		weights[3608] <= 181;
		weights[3609] <= 248;
		weights[3610] <= 98;
		weights[3611] <= 107;
		weights[3612] <= 199;
		weights[3613] <= 198;
		weights[3614] <= 116;
		weights[3615] <= 193;
		weights[3616] <= 220;
		weights[3617] <= 227;
		weights[3618] <= 181;
		weights[3619] <= 234;
		weights[3620] <= 175;
		weights[3621] <= 7;
		weights[3622] <= 19;
		weights[3623] <= 243;
		weights[3624] <= 55;
		weights[3625] <= 127;
		weights[3626] <= 133;
		weights[3627] <= 90;
		weights[3628] <= 129;
		weights[3629] <= 67;
		weights[3630] <= 66;
		weights[3631] <= 17;
		weights[3632] <= 123;
		weights[3633] <= 27;
		weights[3634] <= 28;
		weights[3635] <= 158;
		weights[3636] <= 50;
		weights[3637] <= 146;
		weights[3638] <= 44;
		weights[3639] <= 70;
		weights[3640] <= 194;
		weights[3641] <= 125;
		weights[3642] <= 175;
		weights[3643] <= 242;
		weights[3644] <= 107;
		weights[3645] <= 20;
		weights[3646] <= 125;
		weights[3647] <= 137;
		weights[3648] <= 124;
		weights[3649] <= 212;
		weights[3650] <= 126;
		weights[3651] <= 126;
		weights[3652] <= 106;
		weights[3653] <= 157;
		weights[3654] <= 207;
		weights[3655] <= 110;
		weights[3656] <= 233;
		weights[3657] <= 248;
		weights[3658] <= 14;
		weights[3659] <= 68;
		weights[3660] <= 193;
		weights[3661] <= 244;
		weights[3662] <= 1;
		weights[3663] <= 83;
		weights[3664] <= 223;
		weights[3665] <= 212;
		weights[3666] <= 12;
		weights[3667] <= 183;
		weights[3668] <= 98;
		weights[3669] <= 207;
		weights[3670] <= 102;
		weights[3671] <= 27;
		weights[3672] <= 39;
		weights[3673] <= 127;
		weights[3674] <= 37;
		weights[3675] <= 249;
		weights[3676] <= 237;
		weights[3677] <= 4;
		weights[3678] <= 201;
		weights[3679] <= 20;
		weights[3680] <= 122;
		weights[3681] <= 4;
		weights[3682] <= 73;
		weights[3683] <= 22;
		weights[3684] <= 23;
		weights[3685] <= 250;
		weights[3686] <= 30;
		weights[3687] <= 188;
		weights[3688] <= 181;
		weights[3689] <= 52;
		weights[3690] <= 125;
		weights[3691] <= 238;
		weights[3692] <= 224;
		weights[3693] <= 119;
		weights[3694] <= 35;
		weights[3695] <= 151;
		weights[3696] <= 151;
		weights[3697] <= 222;
		weights[3698] <= 6;
		weights[3699] <= 227;
		weights[3700] <= 235;
		weights[3701] <= 204;
		weights[3702] <= 245;
		weights[3703] <= 232;
		weights[3704] <= 142;
		weights[3705] <= 28;
		weights[3706] <= 143;
		weights[3707] <= 79;
		weights[3708] <= 255;
		weights[3709] <= 236;
		weights[3710] <= 249;
		weights[3711] <= 134;
		weights[3712] <= 129;
		weights[3713] <= 92;
		weights[3714] <= 63;
		weights[3715] <= 188;
		weights[3716] <= 98;
		weights[3717] <= 193;
		weights[3718] <= 54;
		weights[3719] <= 234;
		weights[3720] <= 245;
		weights[3721] <= 95;
		weights[3722] <= 205;
		weights[3723] <= 136;
		weights[3724] <= 67;
		weights[3725] <= 217;
		weights[3726] <= 19;
		weights[3727] <= 151;
		weights[3728] <= 230;
		weights[3729] <= 231;
		weights[3730] <= 122;
		weights[3731] <= 94;
		weights[3732] <= 64;
		weights[3733] <= 200;
		weights[3734] <= 60;
		weights[3735] <= 148;
		weights[3736] <= 128;
		weights[3737] <= 36;
		weights[3738] <= 184;
		weights[3739] <= 166;
		weights[3740] <= 67;
		weights[3741] <= 26;
		weights[3742] <= 150;
		weights[3743] <= 101;
		weights[3744] <= 121;
		weights[3745] <= 246;
		weights[3746] <= 31;
		weights[3747] <= 140;
		weights[3748] <= 6;
		weights[3749] <= 217;
		weights[3750] <= 18;
		weights[3751] <= 69;
		weights[3752] <= 141;
		weights[3753] <= 192;
		weights[3754] <= 140;
		weights[3755] <= 225;
		weights[3756] <= 166;
		weights[3757] <= 227;
		weights[3758] <= 231;
		weights[3759] <= 103;
		weights[3760] <= 8;
		weights[3761] <= 216;
		weights[3762] <= 22;
		weights[3763] <= 13;
		weights[3764] <= 91;
		weights[3765] <= 84;
		weights[3766] <= 160;
		weights[3767] <= 224;
		weights[3768] <= 62;
		weights[3769] <= 151;
		weights[3770] <= 97;
		weights[3771] <= 28;
		weights[3772] <= 145;
		weights[3773] <= 15;
		weights[3774] <= 67;
		weights[3775] <= 43;
		weights[3776] <= 190;
		weights[3777] <= 111;
		weights[3778] <= 51;
		weights[3779] <= 226;
		weights[3780] <= 48;
		weights[3781] <= 144;
		weights[3782] <= 37;
		weights[3783] <= 70;
		weights[3784] <= 153;
		weights[3785] <= 120;
		weights[3786] <= 148;
		weights[3787] <= 47;
		weights[3788] <= 131;
		weights[3789] <= 123;
		weights[3790] <= 228;
		weights[3791] <= 122;
		weights[3792] <= 28;
		weights[3793] <= 146;
		weights[3794] <= 221;
		weights[3795] <= 19;
		weights[3796] <= 6;
		weights[3797] <= 226;
		weights[3798] <= 177;
		weights[3799] <= 13;
		weights[3800] <= 66;
		weights[3801] <= 21;
		weights[3802] <= 182;
		weights[3803] <= 208;
		weights[3804] <= 139;
		weights[3805] <= 135;
		weights[3806] <= 162;
		weights[3807] <= 109;
		weights[3808] <= 251;
		weights[3809] <= 126;
		weights[3810] <= 41;
		weights[3811] <= 23;
		weights[3812] <= 109;
		weights[3813] <= 174;
		weights[3814] <= 125;
		weights[3815] <= 105;
		weights[3816] <= 238;
		weights[3817] <= 222;
		weights[3818] <= 97;
		weights[3819] <= 251;
		weights[3820] <= 162;
		weights[3821] <= 8;
		weights[3822] <= 28;
		weights[3823] <= 208;
		weights[3824] <= 17;
		weights[3825] <= 219;
		weights[3826] <= 111;
		weights[3827] <= 77;
		weights[3828] <= 29;
		weights[3829] <= 78;
		weights[3830] <= 138;
		weights[3831] <= 250;
		weights[3832] <= 62;
		weights[3833] <= 218;
		weights[3834] <= 70;
		weights[3835] <= 213;
		weights[3836] <= 234;
		weights[3837] <= 61;
		weights[3838] <= 171;
		weights[3839] <= 189;
		weights[3840] <= 195;
		weights[3841] <= 42;
		weights[3842] <= 255;
		weights[3843] <= 108;
		weights[3844] <= 101;
		weights[3845] <= 226;
		weights[3846] <= 214;
		weights[3847] <= 225;
		weights[3848] <= 56;
		weights[3849] <= 149;
		weights[3850] <= 171;
		weights[3851] <= 103;
		weights[3852] <= 204;
		weights[3853] <= 69;
		weights[3854] <= 83;
		weights[3855] <= 133;
		weights[3856] <= 105;
		weights[3857] <= 118;
		weights[3858] <= 171;
		weights[3859] <= 230;
		weights[3860] <= 62;
		weights[3861] <= 96;
		weights[3862] <= 200;
		weights[3863] <= 158;
		weights[3864] <= 155;
		weights[3865] <= 196;
		weights[3866] <= 220;
		weights[3867] <= 101;
		weights[3868] <= 89;
		weights[3869] <= 254;
		weights[3870] <= 54;
		weights[3871] <= 148;
		weights[3872] <= 170;
		weights[3873] <= 126;
		weights[3874] <= 106;
		weights[3875] <= 93;
		weights[3876] <= 43;
		weights[3877] <= 60;
		weights[3878] <= 62;
		weights[3879] <= 39;
		weights[3880] <= 103;
		weights[3881] <= 193;
		weights[3882] <= 150;
		weights[3883] <= 12;
		weights[3884] <= 24;
		weights[3885] <= 206;
		weights[3886] <= 217;
		weights[3887] <= 188;
		weights[3888] <= 167;
		weights[3889] <= 6;
		weights[3890] <= 85;
		weights[3891] <= 6;
		weights[3892] <= 82;
		weights[3893] <= 96;
		weights[3894] <= 188;
		weights[3895] <= 111;
		weights[3896] <= 207;
		weights[3897] <= 238;
		weights[3898] <= 63;
		weights[3899] <= 178;
		weights[3900] <= 227;
		weights[3901] <= 23;
		weights[3902] <= 66;
		weights[3903] <= 93;
		weights[3904] <= 63;
		weights[3905] <= 163;
		weights[3906] <= 219;
		weights[3907] <= 187;
		weights[3908] <= 30;
		weights[3909] <= 199;
		weights[3910] <= 41;
		weights[3911] <= 107;
		weights[3912] <= 195;
		weights[3913] <= 162;
		weights[3914] <= 118;
		weights[3915] <= 43;
		weights[3916] <= 14;
		weights[3917] <= 105;
		weights[3918] <= 174;
		weights[3919] <= 146;
		weights[3920] <= 195;
		weights[3921] <= 20;
		weights[3922] <= 6;
		weights[3923] <= 88;
		weights[3924] <= 22;
		weights[3925] <= 144;
		weights[3926] <= 6;
		weights[3927] <= 89;
		weights[3928] <= 163;
		weights[3929] <= 161;
		weights[3930] <= 109;
		weights[3931] <= 104;
		weights[3932] <= 214;
		weights[3933] <= 240;
		weights[3934] <= 240;
		weights[3935] <= 22;
		weights[3936] <= 42;
		weights[3937] <= 179;
		weights[3938] <= 210;
		weights[3939] <= 221;
		weights[3940] <= 148;
		weights[3941] <= 17;
		weights[3942] <= 122;
		weights[3943] <= 4;
		weights[3944] <= 211;
		weights[3945] <= 51;
		weights[3946] <= 69;
		weights[3947] <= 83;
		weights[3948] <= 160;
		weights[3949] <= 28;
		weights[3950] <= 107;
		weights[3951] <= 140;
		weights[3952] <= 236;
		weights[3953] <= 180;
		weights[3954] <= 115;
		weights[3955] <= 56;
		weights[3956] <= 35;
		weights[3957] <= 227;
		weights[3958] <= 143;
		weights[3959] <= 211;
		weights[3960] <= 98;
		weights[3961] <= 55;
		weights[3962] <= 226;
		weights[3963] <= 125;
		weights[3964] <= 186;
		weights[3965] <= 171;
		weights[3966] <= 4;
		weights[3967] <= 123;
		weights[3968] <= 36;
		weights[3969] <= 160;
		weights[3970] <= 17;
		weights[3971] <= 149;
		weights[3972] <= 110;
		weights[3973] <= 246;
		weights[3974] <= 240;
		weights[3975] <= 183;
		weights[3976] <= 6;
		weights[3977] <= 17;
		weights[3978] <= 44;
		weights[3979] <= 252;
		weights[3980] <= 45;
		weights[3981] <= 115;
		weights[3982] <= 120;
		weights[3983] <= 123;
		weights[3984] <= 245;
		weights[3985] <= 124;
		weights[3986] <= 249;
		weights[3987] <= 86;
		weights[3988] <= 106;
		weights[3989] <= 195;
		weights[3990] <= 240;
		weights[3991] <= 255;
		weights[3992] <= 24;
		weights[3993] <= 233;
		weights[3994] <= 70;
		weights[3995] <= 103;
		weights[3996] <= 88;
		weights[3997] <= 130;
		weights[3998] <= 44;
		weights[3999] <= 40;
		weights[4000] <= 196;
		weights[4001] <= 26;
		weights[4002] <= 199;
		weights[4003] <= 123;
		weights[4004] <= 116;
		weights[4005] <= 55;
		weights[4006] <= 24;
		weights[4007] <= 20;
		weights[4008] <= 121;
		weights[4009] <= 58;
		weights[4010] <= 249;
		weights[4011] <= 185;
		weights[4012] <= 247;
		weights[4013] <= 87;
		weights[4014] <= 83;
		weights[4015] <= 8;
		weights[4016] <= 252;
		weights[4017] <= 33;
		weights[4018] <= 129;
		weights[4019] <= 48;
		weights[4020] <= 127;
		weights[4021] <= 181;
		weights[4022] <= 206;
		weights[4023] <= 17;
		weights[4024] <= 25;
		weights[4025] <= 24;
		weights[4026] <= 66;
		weights[4027] <= 91;
		weights[4028] <= 31;
		weights[4029] <= 59;
		weights[4030] <= 33;
		weights[4031] <= 193;
		weights[4032] <= 116;
		weights[4033] <= 66;
		weights[4034] <= 221;
		weights[4035] <= 219;
		weights[4036] <= 109;
		weights[4037] <= 199;
		weights[4038] <= 72;
		weights[4039] <= 198;
		weights[4040] <= 79;
		weights[4041] <= 232;
		weights[4042] <= 108;
		weights[4043] <= 114;
		weights[4044] <= 225;
		weights[4045] <= 85;
		weights[4046] <= 143;
		weights[4047] <= 10;
		weights[4048] <= 46;
		weights[4049] <= 97;
		weights[4050] <= 227;
	end


	always @(negedge(clk)) begin
		if(enable) begin
			case(address)
				12'd0		: data1 <= weights[0];
				12'd1		: data1 <= weights[1];
				12'd2		: data1 <= weights[2];
				12'd3		: data1 <= weights[3];
				12'd4		: data1 <= weights[4];
				12'd5		: data1 <= weights[5];
				12'd6		: data1 <= weights[6];
				12'd7		: data1 <= weights[7];
				12'd8		: data1 <= weights[8];
				12'd9		: data1 <= weights[9];
				12'd10		: data1 <= weights[10];
				12'd11		: data1 <= weights[11];
				12'd12		: data1 <= weights[12];
				12'd13		: data1 <= weights[13];
				12'd14		: data1 <= weights[14];
				12'd15		: data1 <= weights[15];
				12'd16		: data1 <= weights[16];
				12'd17		: data1 <= weights[17];
				12'd18		: data1 <= weights[18];
				12'd19		: data1 <= weights[19];
				12'd20		: data1 <= weights[20];
				12'd21		: data1 <= weights[21];
				12'd22		: data1 <= weights[22];
				12'd23		: data1 <= weights[23];
				12'd24		: data1 <= weights[24];
				12'd25		: data1 <= weights[25];
				12'd26		: data1 <= weights[26];
				12'd27		: data1 <= weights[27];
				12'd28		: data1 <= weights[28];
				12'd29		: data1 <= weights[29];
				12'd30		: data1 <= weights[30];
				12'd31		: data1 <= weights[31];
				12'd32		: data1 <= weights[32];
				12'd33		: data1 <= weights[33];
				12'd34		: data1 <= weights[34];
				12'd35		: data1 <= weights[35];
				12'd36		: data1 <= weights[36];
				12'd37		: data1 <= weights[37];
				12'd38		: data1 <= weights[38];
				12'd39		: data1 <= weights[39];
				12'd40		: data1 <= weights[40];
				12'd41		: data1 <= weights[41];
				12'd42		: data1 <= weights[42];
				12'd43		: data1 <= weights[43];
				12'd44		: data1 <= weights[44];
				12'd45		: data1 <= weights[45];
				12'd46		: data1 <= weights[46];
				12'd47		: data1 <= weights[47];
				12'd48		: data1 <= weights[48];
				12'd49		: data1 <= weights[49];
				12'd50		: data1 <= weights[50];
				12'd51		: data1 <= weights[51];
				12'd52		: data1 <= weights[52];
				12'd53		: data1 <= weights[53];
				12'd54		: data1 <= weights[54];
				12'd55		: data1 <= weights[55];
				12'd56		: data1 <= weights[56];
				12'd57		: data1 <= weights[57];
				12'd58		: data1 <= weights[58];
				12'd59		: data1 <= weights[59];
				12'd60		: data1 <= weights[60];
				12'd61		: data1 <= weights[61];
				12'd62		: data1 <= weights[62];
				12'd63		: data1 <= weights[63];
				12'd64		: data1 <= weights[64];
				12'd65		: data1 <= weights[65];
				12'd66		: data1 <= weights[66];
				12'd67		: data1 <= weights[67];
				12'd68		: data1 <= weights[68];
				12'd69		: data1 <= weights[69];
				12'd70		: data1 <= weights[70];
				12'd71		: data1 <= weights[71];
				12'd72		: data1 <= weights[72];
				12'd73		: data1 <= weights[73];
				12'd74		: data1 <= weights[74];
				12'd75		: data1 <= weights[75];
				12'd76		: data1 <= weights[76];
				12'd77		: data1 <= weights[77];
				12'd78		: data1 <= weights[78];
				12'd79		: data1 <= weights[79];
				12'd80		: data1 <= weights[80];
				12'd81		: data1 <= weights[81];
				12'd82		: data1 <= weights[82];
				12'd83		: data1 <= weights[83];
				12'd84		: data1 <= weights[84];
				12'd85		: data1 <= weights[85];
				12'd86		: data1 <= weights[86];
				12'd87		: data1 <= weights[87];
				12'd88		: data1 <= weights[88];
				12'd89		: data1 <= weights[89];
				12'd90		: data1 <= weights[90];
				12'd91		: data1 <= weights[91];
				12'd92		: data1 <= weights[92];
				12'd93		: data1 <= weights[93];
				12'd94		: data1 <= weights[94];
				12'd95		: data1 <= weights[95];
				12'd96		: data1 <= weights[96];
				12'd97		: data1 <= weights[97];
				12'd98		: data1 <= weights[98];
				12'd99		: data1 <= weights[99];
				12'd100		: data1 <= weights[100];
				12'd101		: data1 <= weights[101];
				12'd102		: data1 <= weights[102];
				12'd103		: data1 <= weights[103];
				12'd104		: data1 <= weights[104];
				12'd105		: data1 <= weights[105];
				12'd106		: data1 <= weights[106];
				12'd107		: data1 <= weights[107];
				12'd108		: data1 <= weights[108];
				12'd109		: data1 <= weights[109];
				12'd110		: data1 <= weights[110];
				12'd111		: data1 <= weights[111];
				12'd112		: data1 <= weights[112];
				12'd113		: data1 <= weights[113];
				12'd114		: data1 <= weights[114];
				12'd115		: data1 <= weights[115];
				12'd116		: data1 <= weights[116];
				12'd117		: data1 <= weights[117];
				12'd118		: data1 <= weights[118];
				12'd119		: data1 <= weights[119];
				12'd120		: data1 <= weights[120];
				12'd121		: data1 <= weights[121];
				12'd122		: data1 <= weights[122];
				12'd123		: data1 <= weights[123];
				12'd124		: data1 <= weights[124];
				12'd125		: data1 <= weights[125];
				12'd126		: data1 <= weights[126];
				12'd127		: data1 <= weights[127];
				12'd128		: data1 <= weights[128];
				12'd129		: data1 <= weights[129];
				12'd130		: data1 <= weights[130];
				12'd131		: data1 <= weights[131];
				12'd132		: data1 <= weights[132];
				12'd133		: data1 <= weights[133];
				12'd134		: data1 <= weights[134];
				12'd135		: data1 <= weights[135];
				12'd136		: data1 <= weights[136];
				12'd137		: data1 <= weights[137];
				12'd138		: data1 <= weights[138];
				12'd139		: data1 <= weights[139];
				12'd140		: data1 <= weights[140];
				12'd141		: data1 <= weights[141];
				12'd142		: data1 <= weights[142];
				12'd143		: data1 <= weights[143];
				12'd144		: data1 <= weights[144];
				12'd145		: data1 <= weights[145];
				12'd146		: data1 <= weights[146];
				12'd147		: data1 <= weights[147];
				12'd148		: data1 <= weights[148];
				12'd149		: data1 <= weights[149];
				12'd150		: data1 <= weights[150];
				12'd151		: data1 <= weights[151];
				12'd152		: data1 <= weights[152];
				12'd153		: data1 <= weights[153];
				12'd154		: data1 <= weights[154];
				12'd155		: data1 <= weights[155];
				12'd156		: data1 <= weights[156];
				12'd157		: data1 <= weights[157];
				12'd158		: data1 <= weights[158];
				12'd159		: data1 <= weights[159];
				12'd160		: data1 <= weights[160];
				12'd161		: data1 <= weights[161];
				12'd162		: data1 <= weights[162];
				12'd163		: data1 <= weights[163];
				12'd164		: data1 <= weights[164];
				12'd165		: data1 <= weights[165];
				12'd166		: data1 <= weights[166];
				12'd167		: data1 <= weights[167];
				12'd168		: data1 <= weights[168];
				12'd169		: data1 <= weights[169];
				12'd170		: data1 <= weights[170];
				12'd171		: data1 <= weights[171];
				12'd172		: data1 <= weights[172];
				12'd173		: data1 <= weights[173];
				12'd174		: data1 <= weights[174];
				12'd175		: data1 <= weights[175];
				12'd176		: data1 <= weights[176];
				12'd177		: data1 <= weights[177];
				12'd178		: data1 <= weights[178];
				12'd179		: data1 <= weights[179];
				12'd180		: data1 <= weights[180];
				12'd181		: data1 <= weights[181];
				12'd182		: data1 <= weights[182];
				12'd183		: data1 <= weights[183];
				12'd184		: data1 <= weights[184];
				12'd185		: data1 <= weights[185];
				12'd186		: data1 <= weights[186];
				12'd187		: data1 <= weights[187];
				12'd188		: data1 <= weights[188];
				12'd189		: data1 <= weights[189];
				12'd190		: data1 <= weights[190];
				12'd191		: data1 <= weights[191];
				12'd192		: data1 <= weights[192];
				12'd193		: data1 <= weights[193];
				12'd194		: data1 <= weights[194];
				12'd195		: data1 <= weights[195];
				12'd196		: data1 <= weights[196];
				12'd197		: data1 <= weights[197];
				12'd198		: data1 <= weights[198];
				12'd199		: data1 <= weights[199];
				12'd200		: data1 <= weights[200];
				12'd201		: data1 <= weights[201];
				12'd202		: data1 <= weights[202];
				12'd203		: data1 <= weights[203];
				12'd204		: data1 <= weights[204];
				12'd205		: data1 <= weights[205];
				12'd206		: data1 <= weights[206];
				12'd207		: data1 <= weights[207];
				12'd208		: data1 <= weights[208];
				12'd209		: data1 <= weights[209];
				12'd210		: data1 <= weights[210];
				12'd211		: data1 <= weights[211];
				12'd212		: data1 <= weights[212];
				12'd213		: data1 <= weights[213];
				12'd214		: data1 <= weights[214];
				12'd215		: data1 <= weights[215];
				12'd216		: data1 <= weights[216];
				12'd217		: data1 <= weights[217];
				12'd218		: data1 <= weights[218];
				12'd219		: data1 <= weights[219];
				12'd220		: data1 <= weights[220];
				12'd221		: data1 <= weights[221];
				12'd222		: data1 <= weights[222];
				12'd223		: data1 <= weights[223];
				12'd224		: data1 <= weights[224];
				12'd225		: data1 <= weights[225];
				12'd226		: data1 <= weights[226];
				12'd227		: data1 <= weights[227];
				12'd228		: data1 <= weights[228];
				12'd229		: data1 <= weights[229];
				12'd230		: data1 <= weights[230];
				12'd231		: data1 <= weights[231];
				12'd232		: data1 <= weights[232];
				12'd233		: data1 <= weights[233];
				12'd234		: data1 <= weights[234];
				12'd235		: data1 <= weights[235];
				12'd236		: data1 <= weights[236];
				12'd237		: data1 <= weights[237];
				12'd238		: data1 <= weights[238];
				12'd239		: data1 <= weights[239];
				12'd240		: data1 <= weights[240];
				12'd241		: data1 <= weights[241];
				12'd242		: data1 <= weights[242];
				12'd243		: data1 <= weights[243];
				12'd244		: data1 <= weights[244];
				12'd245		: data1 <= weights[245];
				12'd246		: data1 <= weights[246];
				12'd247		: data1 <= weights[247];
				12'd248		: data1 <= weights[248];
				12'd249		: data1 <= weights[249];
				12'd250		: data1 <= weights[250];
				12'd251		: data1 <= weights[251];
				12'd252		: data1 <= weights[252];
				12'd253		: data1 <= weights[253];
				12'd254		: data1 <= weights[254];
				12'd255		: data1 <= weights[255];
				12'd256		: data1 <= weights[256];
				12'd257		: data1 <= weights[257];
				12'd258		: data1 <= weights[258];
				12'd259		: data1 <= weights[259];
				12'd260		: data1 <= weights[260];
				12'd261		: data1 <= weights[261];
				12'd262		: data1 <= weights[262];
				12'd263		: data1 <= weights[263];
				12'd264		: data1 <= weights[264];
				12'd265		: data1 <= weights[265];
				12'd266		: data1 <= weights[266];
				12'd267		: data1 <= weights[267];
				12'd268		: data1 <= weights[268];
				12'd269		: data1 <= weights[269];
				12'd270		: data1 <= weights[270];
				12'd271		: data1 <= weights[271];
				12'd272		: data1 <= weights[272];
				12'd273		: data1 <= weights[273];
				12'd274		: data1 <= weights[274];
				12'd275		: data1 <= weights[275];
				12'd276		: data1 <= weights[276];
				12'd277		: data1 <= weights[277];
				12'd278		: data1 <= weights[278];
				12'd279		: data1 <= weights[279];
				12'd280		: data1 <= weights[280];
				12'd281		: data1 <= weights[281];
				12'd282		: data1 <= weights[282];
				12'd283		: data1 <= weights[283];
				12'd284		: data1 <= weights[284];
				12'd285		: data1 <= weights[285];
				12'd286		: data1 <= weights[286];
				12'd287		: data1 <= weights[287];
				12'd288		: data1 <= weights[288];
				12'd289		: data1 <= weights[289];
				12'd290		: data1 <= weights[290];
				12'd291		: data1 <= weights[291];
				12'd292		: data1 <= weights[292];
				12'd293		: data1 <= weights[293];
				12'd294		: data1 <= weights[294];
				12'd295		: data1 <= weights[295];
				12'd296		: data1 <= weights[296];
				12'd297		: data1 <= weights[297];
				12'd298		: data1 <= weights[298];
				12'd299		: data1 <= weights[299];
				12'd300		: data1 <= weights[300];
				12'd301		: data1 <= weights[301];
				12'd302		: data1 <= weights[302];
				12'd303		: data1 <= weights[303];
				12'd304		: data1 <= weights[304];
				12'd305		: data1 <= weights[305];
				12'd306		: data1 <= weights[306];
				12'd307		: data1 <= weights[307];
				12'd308		: data1 <= weights[308];
				12'd309		: data1 <= weights[309];
				12'd310		: data1 <= weights[310];
				12'd311		: data1 <= weights[311];
				12'd312		: data1 <= weights[312];
				12'd313		: data1 <= weights[313];
				12'd314		: data1 <= weights[314];
				12'd315		: data1 <= weights[315];
				12'd316		: data1 <= weights[316];
				12'd317		: data1 <= weights[317];
				12'd318		: data1 <= weights[318];
				12'd319		: data1 <= weights[319];
				12'd320		: data1 <= weights[320];
				12'd321		: data1 <= weights[321];
				12'd322		: data1 <= weights[322];
				12'd323		: data1 <= weights[323];
				12'd324		: data1 <= weights[324];
				12'd325		: data1 <= weights[325];
				12'd326		: data1 <= weights[326];
				12'd327		: data1 <= weights[327];
				12'd328		: data1 <= weights[328];
				12'd329		: data1 <= weights[329];
				12'd330		: data1 <= weights[330];
				12'd331		: data1 <= weights[331];
				12'd332		: data1 <= weights[332];
				12'd333		: data1 <= weights[333];
				12'd334		: data1 <= weights[334];
				12'd335		: data1 <= weights[335];
				12'd336		: data1 <= weights[336];
				12'd337		: data1 <= weights[337];
				12'd338		: data1 <= weights[338];
				12'd339		: data1 <= weights[339];
				12'd340		: data1 <= weights[340];
				12'd341		: data1 <= weights[341];
				12'd342		: data1 <= weights[342];
				12'd343		: data1 <= weights[343];
				12'd344		: data1 <= weights[344];
				12'd345		: data1 <= weights[345];
				12'd346		: data1 <= weights[346];
				12'd347		: data1 <= weights[347];
				12'd348		: data1 <= weights[348];
				12'd349		: data1 <= weights[349];
				12'd350		: data1 <= weights[350];
				12'd351		: data1 <= weights[351];
				12'd352		: data1 <= weights[352];
				12'd353		: data1 <= weights[353];
				12'd354		: data1 <= weights[354];
				12'd355		: data1 <= weights[355];
				12'd356		: data1 <= weights[356];
				12'd357		: data1 <= weights[357];
				12'd358		: data1 <= weights[358];
				12'd359		: data1 <= weights[359];
				12'd360		: data1 <= weights[360];
				12'd361		: data1 <= weights[361];
				12'd362		: data1 <= weights[362];
				12'd363		: data1 <= weights[363];
				12'd364		: data1 <= weights[364];
				12'd365		: data1 <= weights[365];
				12'd366		: data1 <= weights[366];
				12'd367		: data1 <= weights[367];
				12'd368		: data1 <= weights[368];
				12'd369		: data1 <= weights[369];
				12'd370		: data1 <= weights[370];
				12'd371		: data1 <= weights[371];
				12'd372		: data1 <= weights[372];
				12'd373		: data1 <= weights[373];
				12'd374		: data1 <= weights[374];
				12'd375		: data1 <= weights[375];
				12'd376		: data1 <= weights[376];
				12'd377		: data1 <= weights[377];
				12'd378		: data1 <= weights[378];
				12'd379		: data1 <= weights[379];
				12'd380		: data1 <= weights[380];
				12'd381		: data1 <= weights[381];
				12'd382		: data1 <= weights[382];
				12'd383		: data1 <= weights[383];
				12'd384		: data1 <= weights[384];
				12'd385		: data1 <= weights[385];
				12'd386		: data1 <= weights[386];
				12'd387		: data1 <= weights[387];
				12'd388		: data1 <= weights[388];
				12'd389		: data1 <= weights[389];
				12'd390		: data1 <= weights[390];
				12'd391		: data1 <= weights[391];
				12'd392		: data1 <= weights[392];
				12'd393		: data1 <= weights[393];
				12'd394		: data1 <= weights[394];
				12'd395		: data1 <= weights[395];
				12'd396		: data1 <= weights[396];
				12'd397		: data1 <= weights[397];
				12'd398		: data1 <= weights[398];
				12'd399		: data1 <= weights[399];
				12'd400		: data1 <= weights[400];
				12'd401		: data1 <= weights[401];
				12'd402		: data1 <= weights[402];
				12'd403		: data1 <= weights[403];
				12'd404		: data1 <= weights[404];
				12'd405		: data1 <= weights[405];
				12'd406		: data1 <= weights[406];
				12'd407		: data1 <= weights[407];
				12'd408		: data1 <= weights[408];
				12'd409		: data1 <= weights[409];
				12'd410		: data1 <= weights[410];
				12'd411		: data1 <= weights[411];
				12'd412		: data1 <= weights[412];
				12'd413		: data1 <= weights[413];
				12'd414		: data1 <= weights[414];
				12'd415		: data1 <= weights[415];
				12'd416		: data1 <= weights[416];
				12'd417		: data1 <= weights[417];
				12'd418		: data1 <= weights[418];
				12'd419		: data1 <= weights[419];
				12'd420		: data1 <= weights[420];
				12'd421		: data1 <= weights[421];
				12'd422		: data1 <= weights[422];
				12'd423		: data1 <= weights[423];
				12'd424		: data1 <= weights[424];
				12'd425		: data1 <= weights[425];
				12'd426		: data1 <= weights[426];
				12'd427		: data1 <= weights[427];
				12'd428		: data1 <= weights[428];
				12'd429		: data1 <= weights[429];
				12'd430		: data1 <= weights[430];
				12'd431		: data1 <= weights[431];
				12'd432		: data1 <= weights[432];
				12'd433		: data1 <= weights[433];
				12'd434		: data1 <= weights[434];
				12'd435		: data1 <= weights[435];
				12'd436		: data1 <= weights[436];
				12'd437		: data1 <= weights[437];
				12'd438		: data1 <= weights[438];
				12'd439		: data1 <= weights[439];
				12'd440		: data1 <= weights[440];
				12'd441		: data1 <= weights[441];
				12'd442		: data1 <= weights[442];
				12'd443		: data1 <= weights[443];
				12'd444		: data1 <= weights[444];
				12'd445		: data1 <= weights[445];
				12'd446		: data1 <= weights[446];
				12'd447		: data1 <= weights[447];
				12'd448		: data1 <= weights[448];
				12'd449		: data1 <= weights[449];
				12'd450		: data1 <= weights[450];
				12'd451		: data1 <= weights[451];
				12'd452		: data1 <= weights[452];
				12'd453		: data1 <= weights[453];
				12'd454		: data1 <= weights[454];
				12'd455		: data1 <= weights[455];
				12'd456		: data1 <= weights[456];
				12'd457		: data1 <= weights[457];
				12'd458		: data1 <= weights[458];
				12'd459		: data1 <= weights[459];
				12'd460		: data1 <= weights[460];
				12'd461		: data1 <= weights[461];
				12'd462		: data1 <= weights[462];
				12'd463		: data1 <= weights[463];
				12'd464		: data1 <= weights[464];
				12'd465		: data1 <= weights[465];
				12'd466		: data1 <= weights[466];
				12'd467		: data1 <= weights[467];
				12'd468		: data1 <= weights[468];
				12'd469		: data1 <= weights[469];
				12'd470		: data1 <= weights[470];
				12'd471		: data1 <= weights[471];
				12'd472		: data1 <= weights[472];
				12'd473		: data1 <= weights[473];
				12'd474		: data1 <= weights[474];
				12'd475		: data1 <= weights[475];
				12'd476		: data1 <= weights[476];
				12'd477		: data1 <= weights[477];
				12'd478		: data1 <= weights[478];
				12'd479		: data1 <= weights[479];
				12'd480		: data1 <= weights[480];
				12'd481		: data1 <= weights[481];
				12'd482		: data1 <= weights[482];
				12'd483		: data1 <= weights[483];
				12'd484		: data1 <= weights[484];
				12'd485		: data1 <= weights[485];
				12'd486		: data1 <= weights[486];
				12'd487		: data1 <= weights[487];
				12'd488		: data1 <= weights[488];
				12'd489		: data1 <= weights[489];
				12'd490		: data1 <= weights[490];
				12'd491		: data1 <= weights[491];
				12'd492		: data1 <= weights[492];
				12'd493		: data1 <= weights[493];
				12'd494		: data1 <= weights[494];
				12'd495		: data1 <= weights[495];
				12'd496		: data1 <= weights[496];
				12'd497		: data1 <= weights[497];
				12'd498		: data1 <= weights[498];
				12'd499		: data1 <= weights[499];
				12'd500		: data1 <= weights[500];
				12'd501		: data1 <= weights[501];
				12'd502		: data1 <= weights[502];
				12'd503		: data1 <= weights[503];
				12'd504		: data1 <= weights[504];
				12'd505		: data1 <= weights[505];
				12'd506		: data1 <= weights[506];
				12'd507		: data1 <= weights[507];
				12'd508		: data1 <= weights[508];
				12'd509		: data1 <= weights[509];
				12'd510		: data1 <= weights[510];
				12'd511		: data1 <= weights[511];
				12'd512		: data1 <= weights[512];
				12'd513		: data1 <= weights[513];
				12'd514		: data1 <= weights[514];
				12'd515		: data1 <= weights[515];
				12'd516		: data1 <= weights[516];
				12'd517		: data1 <= weights[517];
				12'd518		: data1 <= weights[518];
				12'd519		: data1 <= weights[519];
				12'd520		: data1 <= weights[520];
				12'd521		: data1 <= weights[521];
				12'd522		: data1 <= weights[522];
				12'd523		: data1 <= weights[523];
				12'd524		: data1 <= weights[524];
				12'd525		: data1 <= weights[525];
				12'd526		: data1 <= weights[526];
				12'd527		: data1 <= weights[527];
				12'd528		: data1 <= weights[528];
				12'd529		: data1 <= weights[529];
				12'd530		: data1 <= weights[530];
				12'd531		: data1 <= weights[531];
				12'd532		: data1 <= weights[532];
				12'd533		: data1 <= weights[533];
				12'd534		: data1 <= weights[534];
				12'd535		: data1 <= weights[535];
				12'd536		: data1 <= weights[536];
				12'd537		: data1 <= weights[537];
				12'd538		: data1 <= weights[538];
				12'd539		: data1 <= weights[539];
				12'd540		: data1 <= weights[540];
				12'd541		: data1 <= weights[541];
				12'd542		: data1 <= weights[542];
				12'd543		: data1 <= weights[543];
				12'd544		: data1 <= weights[544];
				12'd545		: data1 <= weights[545];
				12'd546		: data1 <= weights[546];
				12'd547		: data1 <= weights[547];
				12'd548		: data1 <= weights[548];
				12'd549		: data1 <= weights[549];
				12'd550		: data1 <= weights[550];
				12'd551		: data1 <= weights[551];
				12'd552		: data1 <= weights[552];
				12'd553		: data1 <= weights[553];
				12'd554		: data1 <= weights[554];
				12'd555		: data1 <= weights[555];
				12'd556		: data1 <= weights[556];
				12'd557		: data1 <= weights[557];
				12'd558		: data1 <= weights[558];
				12'd559		: data1 <= weights[559];
				12'd560		: data1 <= weights[560];
				12'd561		: data1 <= weights[561];
				12'd562		: data1 <= weights[562];
				12'd563		: data1 <= weights[563];
				12'd564		: data1 <= weights[564];
				12'd565		: data1 <= weights[565];
				12'd566		: data1 <= weights[566];
				12'd567		: data1 <= weights[567];
				12'd568		: data1 <= weights[568];
				12'd569		: data1 <= weights[569];
				12'd570		: data1 <= weights[570];
				12'd571		: data1 <= weights[571];
				12'd572		: data1 <= weights[572];
				12'd573		: data1 <= weights[573];
				12'd574		: data1 <= weights[574];
				12'd575		: data1 <= weights[575];
				12'd576		: data1 <= weights[576];
				12'd577		: data1 <= weights[577];
				12'd578		: data1 <= weights[578];
				12'd579		: data1 <= weights[579];
				12'd580		: data1 <= weights[580];
				12'd581		: data1 <= weights[581];
				12'd582		: data1 <= weights[582];
				12'd583		: data1 <= weights[583];
				12'd584		: data1 <= weights[584];
				12'd585		: data1 <= weights[585];
				12'd586		: data1 <= weights[586];
				12'd587		: data1 <= weights[587];
				12'd588		: data1 <= weights[588];
				12'd589		: data1 <= weights[589];
				12'd590		: data1 <= weights[590];
				12'd591		: data1 <= weights[591];
				12'd592		: data1 <= weights[592];
				12'd593		: data1 <= weights[593];
				12'd594		: data1 <= weights[594];
				12'd595		: data1 <= weights[595];
				12'd596		: data1 <= weights[596];
				12'd597		: data1 <= weights[597];
				12'd598		: data1 <= weights[598];
				12'd599		: data1 <= weights[599];
				12'd600		: data1 <= weights[600];
				12'd601		: data1 <= weights[601];
				12'd602		: data1 <= weights[602];
				12'd603		: data1 <= weights[603];
				12'd604		: data1 <= weights[604];
				12'd605		: data1 <= weights[605];
				12'd606		: data1 <= weights[606];
				12'd607		: data1 <= weights[607];
				12'd608		: data1 <= weights[608];
				12'd609		: data1 <= weights[609];
				12'd610		: data1 <= weights[610];
				12'd611		: data1 <= weights[611];
				12'd612		: data1 <= weights[612];
				12'd613		: data1 <= weights[613];
				12'd614		: data1 <= weights[614];
				12'd615		: data1 <= weights[615];
				12'd616		: data1 <= weights[616];
				12'd617		: data1 <= weights[617];
				12'd618		: data1 <= weights[618];
				12'd619		: data1 <= weights[619];
				12'd620		: data1 <= weights[620];
				12'd621		: data1 <= weights[621];
				12'd622		: data1 <= weights[622];
				12'd623		: data1 <= weights[623];
				12'd624		: data1 <= weights[624];
				12'd625		: data1 <= weights[625];
				12'd626		: data1 <= weights[626];
				12'd627		: data1 <= weights[627];
				12'd628		: data1 <= weights[628];
				12'd629		: data1 <= weights[629];
				12'd630		: data1 <= weights[630];
				12'd631		: data1 <= weights[631];
				12'd632		: data1 <= weights[632];
				12'd633		: data1 <= weights[633];
				12'd634		: data1 <= weights[634];
				12'd635		: data1 <= weights[635];
				12'd636		: data1 <= weights[636];
				12'd637		: data1 <= weights[637];
				12'd638		: data1 <= weights[638];
				12'd639		: data1 <= weights[639];
				12'd640		: data1 <= weights[640];
				12'd641		: data1 <= weights[641];
				12'd642		: data1 <= weights[642];
				12'd643		: data1 <= weights[643];
				12'd644		: data1 <= weights[644];
				12'd645		: data1 <= weights[645];
				12'd646		: data1 <= weights[646];
				12'd647		: data1 <= weights[647];
				12'd648		: data1 <= weights[648];
				12'd649		: data1 <= weights[649];
				12'd650		: data1 <= weights[650];
				12'd651		: data1 <= weights[651];
				12'd652		: data1 <= weights[652];
				12'd653		: data1 <= weights[653];
				12'd654		: data1 <= weights[654];
				12'd655		: data1 <= weights[655];
				12'd656		: data1 <= weights[656];
				12'd657		: data1 <= weights[657];
				12'd658		: data1 <= weights[658];
				12'd659		: data1 <= weights[659];
				12'd660		: data1 <= weights[660];
				12'd661		: data1 <= weights[661];
				12'd662		: data1 <= weights[662];
				12'd663		: data1 <= weights[663];
				12'd664		: data1 <= weights[664];
				12'd665		: data1 <= weights[665];
				12'd666		: data1 <= weights[666];
				12'd667		: data1 <= weights[667];
				12'd668		: data1 <= weights[668];
				12'd669		: data1 <= weights[669];
				12'd670		: data1 <= weights[670];
				12'd671		: data1 <= weights[671];
				12'd672		: data1 <= weights[672];
				12'd673		: data1 <= weights[673];
				12'd674		: data1 <= weights[674];
				12'd675		: data1 <= weights[675];
				12'd676		: data1 <= weights[676];
				12'd677		: data1 <= weights[677];
				12'd678		: data1 <= weights[678];
				12'd679		: data1 <= weights[679];
				12'd680		: data1 <= weights[680];
				12'd681		: data1 <= weights[681];
				12'd682		: data1 <= weights[682];
				12'd683		: data1 <= weights[683];
				12'd684		: data1 <= weights[684];
				12'd685		: data1 <= weights[685];
				12'd686		: data1 <= weights[686];
				12'd687		: data1 <= weights[687];
				12'd688		: data1 <= weights[688];
				12'd689		: data1 <= weights[689];
				12'd690		: data1 <= weights[690];
				12'd691		: data1 <= weights[691];
				12'd692		: data1 <= weights[692];
				12'd693		: data1 <= weights[693];
				12'd694		: data1 <= weights[694];
				12'd695		: data1 <= weights[695];
				12'd696		: data1 <= weights[696];
				12'd697		: data1 <= weights[697];
				12'd698		: data1 <= weights[698];
				12'd699		: data1 <= weights[699];
				12'd700		: data1 <= weights[700];
				12'd701		: data1 <= weights[701];
				12'd702		: data1 <= weights[702];
				12'd703		: data1 <= weights[703];
				12'd704		: data1 <= weights[704];
				12'd705		: data1 <= weights[705];
				12'd706		: data1 <= weights[706];
				12'd707		: data1 <= weights[707];
				12'd708		: data1 <= weights[708];
				12'd709		: data1 <= weights[709];
				12'd710		: data1 <= weights[710];
				12'd711		: data1 <= weights[711];
				12'd712		: data1 <= weights[712];
				12'd713		: data1 <= weights[713];
				12'd714		: data1 <= weights[714];
				12'd715		: data1 <= weights[715];
				12'd716		: data1 <= weights[716];
				12'd717		: data1 <= weights[717];
				12'd718		: data1 <= weights[718];
				12'd719		: data1 <= weights[719];
				12'd720		: data1 <= weights[720];
				12'd721		: data1 <= weights[721];
				12'd722		: data1 <= weights[722];
				12'd723		: data1 <= weights[723];
				12'd724		: data1 <= weights[724];
				12'd725		: data1 <= weights[725];
				12'd726		: data1 <= weights[726];
				12'd727		: data1 <= weights[727];
				12'd728		: data1 <= weights[728];
				12'd729		: data1 <= weights[729];
				12'd730		: data1 <= weights[730];
				12'd731		: data1 <= weights[731];
				12'd732		: data1 <= weights[732];
				12'd733		: data1 <= weights[733];
				12'd734		: data1 <= weights[734];
				12'd735		: data1 <= weights[735];
				12'd736		: data1 <= weights[736];
				12'd737		: data1 <= weights[737];
				12'd738		: data1 <= weights[738];
				12'd739		: data1 <= weights[739];
				12'd740		: data1 <= weights[740];
				12'd741		: data1 <= weights[741];
				12'd742		: data1 <= weights[742];
				12'd743		: data1 <= weights[743];
				12'd744		: data1 <= weights[744];
				12'd745		: data1 <= weights[745];
				12'd746		: data1 <= weights[746];
				12'd747		: data1 <= weights[747];
				12'd748		: data1 <= weights[748];
				12'd749		: data1 <= weights[749];
				12'd750		: data1 <= weights[750];
				12'd751		: data1 <= weights[751];
				12'd752		: data1 <= weights[752];
				12'd753		: data1 <= weights[753];
				12'd754		: data1 <= weights[754];
				12'd755		: data1 <= weights[755];
				12'd756		: data1 <= weights[756];
				12'd757		: data1 <= weights[757];
				12'd758		: data1 <= weights[758];
				12'd759		: data1 <= weights[759];
				12'd760		: data1 <= weights[760];
				12'd761		: data1 <= weights[761];
				12'd762		: data1 <= weights[762];
				12'd763		: data1 <= weights[763];
				12'd764		: data1 <= weights[764];
				12'd765		: data1 <= weights[765];
				12'd766		: data1 <= weights[766];
				12'd767		: data1 <= weights[767];
				12'd768		: data1 <= weights[768];
				12'd769		: data1 <= weights[769];
				12'd770		: data1 <= weights[770];
				12'd771		: data1 <= weights[771];
				12'd772		: data1 <= weights[772];
				12'd773		: data1 <= weights[773];
				12'd774		: data1 <= weights[774];
				12'd775		: data1 <= weights[775];
				12'd776		: data1 <= weights[776];
				12'd777		: data1 <= weights[777];
				12'd778		: data1 <= weights[778];
				12'd779		: data1 <= weights[779];
				12'd780		: data1 <= weights[780];
				12'd781		: data1 <= weights[781];
				12'd782		: data1 <= weights[782];
				12'd783		: data1 <= weights[783];
				12'd784		: data1 <= weights[784];
				12'd785		: data1 <= weights[785];
				12'd786		: data1 <= weights[786];
				12'd787		: data1 <= weights[787];
				12'd788		: data1 <= weights[788];
				12'd789		: data1 <= weights[789];
				12'd790		: data1 <= weights[790];
				12'd791		: data1 <= weights[791];
				12'd792		: data1 <= weights[792];
				12'd793		: data1 <= weights[793];
				12'd794		: data1 <= weights[794];
				12'd795		: data1 <= weights[795];
				12'd796		: data1 <= weights[796];
				12'd797		: data1 <= weights[797];
				12'd798		: data1 <= weights[798];
				12'd799		: data1 <= weights[799];
				12'd800		: data1 <= weights[800];
				12'd801		: data1 <= weights[801];
				12'd802		: data1 <= weights[802];
				12'd803		: data1 <= weights[803];
				12'd804		: data1 <= weights[804];
				12'd805		: data1 <= weights[805];
				12'd806		: data1 <= weights[806];
				12'd807		: data1 <= weights[807];
				12'd808		: data1 <= weights[808];
				12'd809		: data1 <= weights[809];
				12'd810		: data1 <= weights[810];
				12'd811		: data1 <= weights[811];
				12'd812		: data1 <= weights[812];
				12'd813		: data1 <= weights[813];
				12'd814		: data1 <= weights[814];
				12'd815		: data1 <= weights[815];
				12'd816		: data1 <= weights[816];
				12'd817		: data1 <= weights[817];
				12'd818		: data1 <= weights[818];
				12'd819		: data1 <= weights[819];
				12'd820		: data1 <= weights[820];
				12'd821		: data1 <= weights[821];
				12'd822		: data1 <= weights[822];
				12'd823		: data1 <= weights[823];
				12'd824		: data1 <= weights[824];
				12'd825		: data1 <= weights[825];
				12'd826		: data1 <= weights[826];
				12'd827		: data1 <= weights[827];
				12'd828		: data1 <= weights[828];
				12'd829		: data1 <= weights[829];
				12'd830		: data1 <= weights[830];
				12'd831		: data1 <= weights[831];
				12'd832		: data1 <= weights[832];
				12'd833		: data1 <= weights[833];
				12'd834		: data1 <= weights[834];
				12'd835		: data1 <= weights[835];
				12'd836		: data1 <= weights[836];
				12'd837		: data1 <= weights[837];
				12'd838		: data1 <= weights[838];
				12'd839		: data1 <= weights[839];
				12'd840		: data1 <= weights[840];
				12'd841		: data1 <= weights[841];
				12'd842		: data1 <= weights[842];
				12'd843		: data1 <= weights[843];
				12'd844		: data1 <= weights[844];
				12'd845		: data1 <= weights[845];
				12'd846		: data1 <= weights[846];
				12'd847		: data1 <= weights[847];
				12'd848		: data1 <= weights[848];
				12'd849		: data1 <= weights[849];
				12'd850		: data1 <= weights[850];
				12'd851		: data1 <= weights[851];
				12'd852		: data1 <= weights[852];
				12'd853		: data1 <= weights[853];
				12'd854		: data1 <= weights[854];
				12'd855		: data1 <= weights[855];
				12'd856		: data1 <= weights[856];
				12'd857		: data1 <= weights[857];
				12'd858		: data1 <= weights[858];
				12'd859		: data1 <= weights[859];
				12'd860		: data1 <= weights[860];
				12'd861		: data1 <= weights[861];
				12'd862		: data1 <= weights[862];
				12'd863		: data1 <= weights[863];
				12'd864		: data1 <= weights[864];
				12'd865		: data1 <= weights[865];
				12'd866		: data1 <= weights[866];
				12'd867		: data1 <= weights[867];
				12'd868		: data1 <= weights[868];
				12'd869		: data1 <= weights[869];
				12'd870		: data1 <= weights[870];
				12'd871		: data1 <= weights[871];
				12'd872		: data1 <= weights[872];
				12'd873		: data1 <= weights[873];
				12'd874		: data1 <= weights[874];
				12'd875		: data1 <= weights[875];
				12'd876		: data1 <= weights[876];
				12'd877		: data1 <= weights[877];
				12'd878		: data1 <= weights[878];
				12'd879		: data1 <= weights[879];
				12'd880		: data1 <= weights[880];
				12'd881		: data1 <= weights[881];
				12'd882		: data1 <= weights[882];
				12'd883		: data1 <= weights[883];
				12'd884		: data1 <= weights[884];
				12'd885		: data1 <= weights[885];
				12'd886		: data1 <= weights[886];
				12'd887		: data1 <= weights[887];
				12'd888		: data1 <= weights[888];
				12'd889		: data1 <= weights[889];
				12'd890		: data1 <= weights[890];
				12'd891		: data1 <= weights[891];
				12'd892		: data1 <= weights[892];
				12'd893		: data1 <= weights[893];
				12'd894		: data1 <= weights[894];
				12'd895		: data1 <= weights[895];
				12'd896		: data1 <= weights[896];
				12'd897		: data1 <= weights[897];
				12'd898		: data1 <= weights[898];
				12'd899		: data1 <= weights[899];
				12'd900		: data1 <= weights[900];
				12'd901		: data1 <= weights[901];
				12'd902		: data1 <= weights[902];
				12'd903		: data1 <= weights[903];
				12'd904		: data1 <= weights[904];
				12'd905		: data1 <= weights[905];
				12'd906		: data1 <= weights[906];
				12'd907		: data1 <= weights[907];
				12'd908		: data1 <= weights[908];
				12'd909		: data1 <= weights[909];
				12'd910		: data1 <= weights[910];
				12'd911		: data1 <= weights[911];
				12'd912		: data1 <= weights[912];
				12'd913		: data1 <= weights[913];
				12'd914		: data1 <= weights[914];
				12'd915		: data1 <= weights[915];
				12'd916		: data1 <= weights[916];
				12'd917		: data1 <= weights[917];
				12'd918		: data1 <= weights[918];
				12'd919		: data1 <= weights[919];
				12'd920		: data1 <= weights[920];
				12'd921		: data1 <= weights[921];
				12'd922		: data1 <= weights[922];
				12'd923		: data1 <= weights[923];
				12'd924		: data1 <= weights[924];
				12'd925		: data1 <= weights[925];
				12'd926		: data1 <= weights[926];
				12'd927		: data1 <= weights[927];
				12'd928		: data1 <= weights[928];
				12'd929		: data1 <= weights[929];
				12'd930		: data1 <= weights[930];
				12'd931		: data1 <= weights[931];
				12'd932		: data1 <= weights[932];
				12'd933		: data1 <= weights[933];
				12'd934		: data1 <= weights[934];
				12'd935		: data1 <= weights[935];
				12'd936		: data1 <= weights[936];
				12'd937		: data1 <= weights[937];
				12'd938		: data1 <= weights[938];
				12'd939		: data1 <= weights[939];
				12'd940		: data1 <= weights[940];
				12'd941		: data1 <= weights[941];
				12'd942		: data1 <= weights[942];
				12'd943		: data1 <= weights[943];
				12'd944		: data1 <= weights[944];
				12'd945		: data1 <= weights[945];
				12'd946		: data1 <= weights[946];
				12'd947		: data1 <= weights[947];
				12'd948		: data1 <= weights[948];
				12'd949		: data1 <= weights[949];
				12'd950		: data1 <= weights[950];
				12'd951		: data1 <= weights[951];
				12'd952		: data1 <= weights[952];
				12'd953		: data1 <= weights[953];
				12'd954		: data1 <= weights[954];
				12'd955		: data1 <= weights[955];
				12'd956		: data1 <= weights[956];
				12'd957		: data1 <= weights[957];
				12'd958		: data1 <= weights[958];
				12'd959		: data1 <= weights[959];
				12'd960		: data1 <= weights[960];
				12'd961		: data1 <= weights[961];
				12'd962		: data1 <= weights[962];
				12'd963		: data1 <= weights[963];
				12'd964		: data1 <= weights[964];
				12'd965		: data1 <= weights[965];
				12'd966		: data1 <= weights[966];
				12'd967		: data1 <= weights[967];
				12'd968		: data1 <= weights[968];
				12'd969		: data1 <= weights[969];
				12'd970		: data1 <= weights[970];
				12'd971		: data1 <= weights[971];
				12'd972		: data1 <= weights[972];
				12'd973		: data1 <= weights[973];
				12'd974		: data1 <= weights[974];
				12'd975		: data1 <= weights[975];
				12'd976		: data1 <= weights[976];
				12'd977		: data1 <= weights[977];
				12'd978		: data1 <= weights[978];
				12'd979		: data1 <= weights[979];
				12'd980		: data1 <= weights[980];
				12'd981		: data1 <= weights[981];
				12'd982		: data1 <= weights[982];
				12'd983		: data1 <= weights[983];
				12'd984		: data1 <= weights[984];
				12'd985		: data1 <= weights[985];
				12'd986		: data1 <= weights[986];
				12'd987		: data1 <= weights[987];
				12'd988		: data1 <= weights[988];
				12'd989		: data1 <= weights[989];
				12'd990		: data1 <= weights[990];
				12'd991		: data1 <= weights[991];
				12'd992		: data1 <= weights[992];
				12'd993		: data1 <= weights[993];
				12'd994		: data1 <= weights[994];
				12'd995		: data1 <= weights[995];
				12'd996		: data1 <= weights[996];
				12'd997		: data1 <= weights[997];
				12'd998		: data1 <= weights[998];
				12'd999		: data1 <= weights[999];
				12'd1000	: data1 <= weights[1000];
				12'd1001	: data1 <= weights[1001];
				12'd1002	: data1 <= weights[1002];
				12'd1003	: data1 <= weights[1003];
				12'd1004	: data1 <= weights[1004];
				12'd1005	: data1 <= weights[1005];
				12'd1006	: data1 <= weights[1006];
				12'd1007	: data1 <= weights[1007];
				12'd1008	: data1 <= weights[1008];
				12'd1009	: data1 <= weights[1009];
				12'd1010	: data1 <= weights[1010];
				12'd1011	: data1 <= weights[1011];
				12'd1012	: data1 <= weights[1012];
				12'd1013	: data1 <= weights[1013];
				12'd1014	: data1 <= weights[1014];
				12'd1015	: data1 <= weights[1015];
				12'd1016	: data1 <= weights[1016];
				12'd1017	: data1 <= weights[1017];
				12'd1018	: data1 <= weights[1018];
				12'd1019	: data1 <= weights[1019];
				12'd1020	: data1 <= weights[1020];
				12'd1021	: data1 <= weights[1021];
				12'd1022	: data1 <= weights[1022];
				12'd1023	: data1 <= weights[1023];
				12'd1024	: data1 <= weights[1024];
				12'd1025	: data1 <= weights[1025];
				12'd1026	: data1 <= weights[1026];
				12'd1027	: data1 <= weights[1027];
				12'd1028	: data1 <= weights[1028];
				12'd1029	: data1 <= weights[1029];
				12'd1030	: data1 <= weights[1030];
				12'd1031	: data1 <= weights[1031];
				12'd1032	: data1 <= weights[1032];
				12'd1033	: data1 <= weights[1033];
				12'd1034	: data1 <= weights[1034];
				12'd1035	: data1 <= weights[1035];
				12'd1036	: data1 <= weights[1036];
				12'd1037	: data1 <= weights[1037];
				12'd1038	: data1 <= weights[1038];
				12'd1039	: data1 <= weights[1039];
				12'd1040	: data1 <= weights[1040];
				12'd1041	: data1 <= weights[1041];
				12'd1042	: data1 <= weights[1042];
				12'd1043	: data1 <= weights[1043];
				12'd1044	: data1 <= weights[1044];
				12'd1045	: data1 <= weights[1045];
				12'd1046	: data1 <= weights[1046];
				12'd1047	: data1 <= weights[1047];
				12'd1048	: data1 <= weights[1048];
				12'd1049	: data1 <= weights[1049];
				12'd1050	: data1 <= weights[1050];
				12'd1051	: data1 <= weights[1051];
				12'd1052	: data1 <= weights[1052];
				12'd1053	: data1 <= weights[1053];
				12'd1054	: data1 <= weights[1054];
				12'd1055	: data1 <= weights[1055];
				12'd1056	: data1 <= weights[1056];
				12'd1057	: data1 <= weights[1057];
				12'd1058	: data1 <= weights[1058];
				12'd1059	: data1 <= weights[1059];
				12'd1060	: data1 <= weights[1060];
				12'd1061	: data1 <= weights[1061];
				12'd1062	: data1 <= weights[1062];
				12'd1063	: data1 <= weights[1063];
				12'd1064	: data1 <= weights[1064];
				12'd1065	: data1 <= weights[1065];
				12'd1066	: data1 <= weights[1066];
				12'd1067	: data1 <= weights[1067];
				12'd1068	: data1 <= weights[1068];
				12'd1069	: data1 <= weights[1069];
				12'd1070	: data1 <= weights[1070];
				12'd1071	: data1 <= weights[1071];
				12'd1072	: data1 <= weights[1072];
				12'd1073	: data1 <= weights[1073];
				12'd1074	: data1 <= weights[1074];
				12'd1075	: data1 <= weights[1075];
				12'd1076	: data1 <= weights[1076];
				12'd1077	: data1 <= weights[1077];
				12'd1078	: data1 <= weights[1078];
				12'd1079	: data1 <= weights[1079];
				12'd1080	: data1 <= weights[1080];
				12'd1081	: data1 <= weights[1081];
				12'd1082	: data1 <= weights[1082];
				12'd1083	: data1 <= weights[1083];
				12'd1084	: data1 <= weights[1084];
				12'd1085	: data1 <= weights[1085];
				12'd1086	: data1 <= weights[1086];
				12'd1087	: data1 <= weights[1087];
				12'd1088	: data1 <= weights[1088];
				12'd1089	: data1 <= weights[1089];
				12'd1090	: data1 <= weights[1090];
				12'd1091	: data1 <= weights[1091];
				12'd1092	: data1 <= weights[1092];
				12'd1093	: data1 <= weights[1093];
				12'd1094	: data1 <= weights[1094];
				12'd1095	: data1 <= weights[1095];
				12'd1096	: data1 <= weights[1096];
				12'd1097	: data1 <= weights[1097];
				12'd1098	: data1 <= weights[1098];
				12'd1099	: data1 <= weights[1099];
				12'd1100	: data1 <= weights[1100];
				12'd1101	: data1 <= weights[1101];
				12'd1102	: data1 <= weights[1102];
				12'd1103	: data1 <= weights[1103];
				12'd1104	: data1 <= weights[1104];
				12'd1105	: data1 <= weights[1105];
				12'd1106	: data1 <= weights[1106];
				12'd1107	: data1 <= weights[1107];
				12'd1108	: data1 <= weights[1108];
				12'd1109	: data1 <= weights[1109];
				12'd1110	: data1 <= weights[1110];
				12'd1111	: data1 <= weights[1111];
				12'd1112	: data1 <= weights[1112];
				12'd1113	: data1 <= weights[1113];
				12'd1114	: data1 <= weights[1114];
				12'd1115	: data1 <= weights[1115];
				12'd1116	: data1 <= weights[1116];
				12'd1117	: data1 <= weights[1117];
				12'd1118	: data1 <= weights[1118];
				12'd1119	: data1 <= weights[1119];
				12'd1120	: data1 <= weights[1120];
				12'd1121	: data1 <= weights[1121];
				12'd1122	: data1 <= weights[1122];
				12'd1123	: data1 <= weights[1123];
				12'd1124	: data1 <= weights[1124];
				12'd1125	: data1 <= weights[1125];
				12'd1126	: data1 <= weights[1126];
				12'd1127	: data1 <= weights[1127];
				12'd1128	: data1 <= weights[1128];
				12'd1129	: data1 <= weights[1129];
				12'd1130	: data1 <= weights[1130];
				12'd1131	: data1 <= weights[1131];
				12'd1132	: data1 <= weights[1132];
				12'd1133	: data1 <= weights[1133];
				12'd1134	: data1 <= weights[1134];
				12'd1135	: data1 <= weights[1135];
				12'd1136	: data1 <= weights[1136];
				12'd1137	: data1 <= weights[1137];
				12'd1138	: data1 <= weights[1138];
				12'd1139	: data1 <= weights[1139];
				12'd1140	: data1 <= weights[1140];
				12'd1141	: data1 <= weights[1141];
				12'd1142	: data1 <= weights[1142];
				12'd1143	: data1 <= weights[1143];
				12'd1144	: data1 <= weights[1144];
				12'd1145	: data1 <= weights[1145];
				12'd1146	: data1 <= weights[1146];
				12'd1147	: data1 <= weights[1147];
				12'd1148	: data1 <= weights[1148];
				12'd1149	: data1 <= weights[1149];
				12'd1150	: data1 <= weights[1150];
				12'd1151	: data1 <= weights[1151];
				12'd1152	: data1 <= weights[1152];
				12'd1153	: data1 <= weights[1153];
				12'd1154	: data1 <= weights[1154];
				12'd1155	: data1 <= weights[1155];
				12'd1156	: data1 <= weights[1156];
				12'd1157	: data1 <= weights[1157];
				12'd1158	: data1 <= weights[1158];
				12'd1159	: data1 <= weights[1159];
				12'd1160	: data1 <= weights[1160];
				12'd1161	: data1 <= weights[1161];
				12'd1162	: data1 <= weights[1162];
				12'd1163	: data1 <= weights[1163];
				12'd1164	: data1 <= weights[1164];
				12'd1165	: data1 <= weights[1165];
				12'd1166	: data1 <= weights[1166];
				12'd1167	: data1 <= weights[1167];
				12'd1168	: data1 <= weights[1168];
				12'd1169	: data1 <= weights[1169];
				12'd1170	: data1 <= weights[1170];
				12'd1171	: data1 <= weights[1171];
				12'd1172	: data1 <= weights[1172];
				12'd1173	: data1 <= weights[1173];
				12'd1174	: data1 <= weights[1174];
				12'd1175	: data1 <= weights[1175];
				12'd1176	: data1 <= weights[1176];
				12'd1177	: data1 <= weights[1177];
				12'd1178	: data1 <= weights[1178];
				12'd1179	: data1 <= weights[1179];
				12'd1180	: data1 <= weights[1180];
				12'd1181	: data1 <= weights[1181];
				12'd1182	: data1 <= weights[1182];
				12'd1183	: data1 <= weights[1183];
				12'd1184	: data1 <= weights[1184];
				12'd1185	: data1 <= weights[1185];
				12'd1186	: data1 <= weights[1186];
				12'd1187	: data1 <= weights[1187];
				12'd1188	: data1 <= weights[1188];
				12'd1189	: data1 <= weights[1189];
				12'd1190	: data1 <= weights[1190];
				12'd1191	: data1 <= weights[1191];
				12'd1192	: data1 <= weights[1192];
				12'd1193	: data1 <= weights[1193];
				12'd1194	: data1 <= weights[1194];
				12'd1195	: data1 <= weights[1195];
				12'd1196	: data1 <= weights[1196];
				12'd1197	: data1 <= weights[1197];
				12'd1198	: data1 <= weights[1198];
				12'd1199	: data1 <= weights[1199];
				12'd1200	: data1 <= weights[1200];
				12'd1201	: data1 <= weights[1201];
				12'd1202	: data1 <= weights[1202];
				12'd1203	: data1 <= weights[1203];
				12'd1204	: data1 <= weights[1204];
				12'd1205	: data1 <= weights[1205];
				12'd1206	: data1 <= weights[1206];
				12'd1207	: data1 <= weights[1207];
				12'd1208	: data1 <= weights[1208];
				12'd1209	: data1 <= weights[1209];
				12'd1210	: data1 <= weights[1210];
				12'd1211	: data1 <= weights[1211];
				12'd1212	: data1 <= weights[1212];
				12'd1213	: data1 <= weights[1213];
				12'd1214	: data1 <= weights[1214];
				12'd1215	: data1 <= weights[1215];
				12'd1216	: data1 <= weights[1216];
				12'd1217	: data1 <= weights[1217];
				12'd1218	: data1 <= weights[1218];
				12'd1219	: data1 <= weights[1219];
				12'd1220	: data1 <= weights[1220];
				12'd1221	: data1 <= weights[1221];
				12'd1222	: data1 <= weights[1222];
				12'd1223	: data1 <= weights[1223];
				12'd1224	: data1 <= weights[1224];
				12'd1225	: data1 <= weights[1225];
				12'd1226	: data1 <= weights[1226];
				12'd1227	: data1 <= weights[1227];
				12'd1228	: data1 <= weights[1228];
				12'd1229	: data1 <= weights[1229];
				12'd1230	: data1 <= weights[1230];
				12'd1231	: data1 <= weights[1231];
				12'd1232	: data1 <= weights[1232];
				12'd1233	: data1 <= weights[1233];
				12'd1234	: data1 <= weights[1234];
				12'd1235	: data1 <= weights[1235];
				12'd1236	: data1 <= weights[1236];
				12'd1237	: data1 <= weights[1237];
				12'd1238	: data1 <= weights[1238];
				12'd1239	: data1 <= weights[1239];
				12'd1240	: data1 <= weights[1240];
				12'd1241	: data1 <= weights[1241];
				12'd1242	: data1 <= weights[1242];
				12'd1243	: data1 <= weights[1243];
				12'd1244	: data1 <= weights[1244];
				12'd1245	: data1 <= weights[1245];
				12'd1246	: data1 <= weights[1246];
				12'd1247	: data1 <= weights[1247];
				12'd1248	: data1 <= weights[1248];
				12'd1249	: data1 <= weights[1249];
				12'd1250	: data1 <= weights[1250];
				12'd1251	: data1 <= weights[1251];
				12'd1252	: data1 <= weights[1252];
				12'd1253	: data1 <= weights[1253];
				12'd1254	: data1 <= weights[1254];
				12'd1255	: data1 <= weights[1255];
				12'd1256	: data1 <= weights[1256];
				12'd1257	: data1 <= weights[1257];
				12'd1258	: data1 <= weights[1258];
				12'd1259	: data1 <= weights[1259];
				12'd1260	: data1 <= weights[1260];
				12'd1261	: data1 <= weights[1261];
				12'd1262	: data1 <= weights[1262];
				12'd1263	: data1 <= weights[1263];
				12'd1264	: data1 <= weights[1264];
				12'd1265	: data1 <= weights[1265];
				12'd1266	: data1 <= weights[1266];
				12'd1267	: data1 <= weights[1267];
				12'd1268	: data1 <= weights[1268];
				12'd1269	: data1 <= weights[1269];
				12'd1270	: data1 <= weights[1270];
				12'd1271	: data1 <= weights[1271];
				12'd1272	: data1 <= weights[1272];
				12'd1273	: data1 <= weights[1273];
				12'd1274	: data1 <= weights[1274];
				12'd1275	: data1 <= weights[1275];
				12'd1276	: data1 <= weights[1276];
				12'd1277	: data1 <= weights[1277];
				12'd1278	: data1 <= weights[1278];
				12'd1279	: data1 <= weights[1279];
				12'd1280	: data1 <= weights[1280];
				12'd1281	: data1 <= weights[1281];
				12'd1282	: data1 <= weights[1282];
				12'd1283	: data1 <= weights[1283];
				12'd1284	: data1 <= weights[1284];
				12'd1285	: data1 <= weights[1285];
				12'd1286	: data1 <= weights[1286];
				12'd1287	: data1 <= weights[1287];
				12'd1288	: data1 <= weights[1288];
				12'd1289	: data1 <= weights[1289];
				12'd1290	: data1 <= weights[1290];
				12'd1291	: data1 <= weights[1291];
				12'd1292	: data1 <= weights[1292];
				12'd1293	: data1 <= weights[1293];
				12'd1294	: data1 <= weights[1294];
				12'd1295	: data1 <= weights[1295];
				12'd1296	: data1 <= weights[1296];
				12'd1297	: data1 <= weights[1297];
				12'd1298	: data1 <= weights[1298];
				12'd1299	: data1 <= weights[1299];
				12'd1300	: data1 <= weights[1300];
				12'd1301	: data1 <= weights[1301];
				12'd1302	: data1 <= weights[1302];
				12'd1303	: data1 <= weights[1303];
				12'd1304	: data1 <= weights[1304];
				12'd1305	: data1 <= weights[1305];
				12'd1306	: data1 <= weights[1306];
				12'd1307	: data1 <= weights[1307];
				12'd1308	: data1 <= weights[1308];
				12'd1309	: data1 <= weights[1309];
				12'd1310	: data1 <= weights[1310];
				12'd1311	: data1 <= weights[1311];
				12'd1312	: data1 <= weights[1312];
				12'd1313	: data1 <= weights[1313];
				12'd1314	: data1 <= weights[1314];
				12'd1315	: data1 <= weights[1315];
				12'd1316	: data1 <= weights[1316];
				12'd1317	: data1 <= weights[1317];
				12'd1318	: data1 <= weights[1318];
				12'd1319	: data1 <= weights[1319];
				12'd1320	: data1 <= weights[1320];
				12'd1321	: data1 <= weights[1321];
				12'd1322	: data1 <= weights[1322];
				12'd1323	: data1 <= weights[1323];
				12'd1324	: data1 <= weights[1324];
				12'd1325	: data1 <= weights[1325];
				12'd1326	: data1 <= weights[1326];
				12'd1327	: data1 <= weights[1327];
				12'd1328	: data1 <= weights[1328];
				12'd1329	: data1 <= weights[1329];
				12'd1330	: data1 <= weights[1330];
				12'd1331	: data1 <= weights[1331];
				12'd1332	: data1 <= weights[1332];
				12'd1333	: data1 <= weights[1333];
				12'd1334	: data1 <= weights[1334];
				12'd1335	: data1 <= weights[1335];
				12'd1336	: data1 <= weights[1336];
				12'd1337	: data1 <= weights[1337];
				12'd1338	: data1 <= weights[1338];
				12'd1339	: data1 <= weights[1339];
				12'd1340	: data1 <= weights[1340];
				12'd1341	: data1 <= weights[1341];
				12'd1342	: data1 <= weights[1342];
				12'd1343	: data1 <= weights[1343];
				12'd1344	: data1 <= weights[1344];
				12'd1345	: data1 <= weights[1345];
				12'd1346	: data1 <= weights[1346];
				12'd1347	: data1 <= weights[1347];
				12'd1348	: data1 <= weights[1348];
				12'd1349	: data1 <= weights[1349];
				12'd1350	: data1 <= weights[1350];
				12'd1351	: data1 <= weights[1351];
				12'd1352	: data1 <= weights[1352];
				12'd1353	: data1 <= weights[1353];
				12'd1354	: data1 <= weights[1354];
				12'd1355	: data1 <= weights[1355];
				12'd1356	: data1 <= weights[1356];
				12'd1357	: data1 <= weights[1357];
				12'd1358	: data1 <= weights[1358];
				12'd1359	: data1 <= weights[1359];
				12'd1360	: data1 <= weights[1360];
				12'd1361	: data1 <= weights[1361];
				12'd1362	: data1 <= weights[1362];
				12'd1363	: data1 <= weights[1363];
				12'd1364	: data1 <= weights[1364];
				12'd1365	: data1 <= weights[1365];
				12'd1366	: data1 <= weights[1366];
				12'd1367	: data1 <= weights[1367];
				12'd1368	: data1 <= weights[1368];
				12'd1369	: data1 <= weights[1369];
				12'd1370	: data1 <= weights[1370];
				12'd1371	: data1 <= weights[1371];
				12'd1372	: data1 <= weights[1372];
				12'd1373	: data1 <= weights[1373];
				12'd1374	: data1 <= weights[1374];
				12'd1375	: data1 <= weights[1375];
				12'd1376	: data1 <= weights[1376];
				12'd1377	: data1 <= weights[1377];
				12'd1378	: data1 <= weights[1378];
				12'd1379	: data1 <= weights[1379];
				12'd1380	: data1 <= weights[1380];
				12'd1381	: data1 <= weights[1381];
				12'd1382	: data1 <= weights[1382];
				12'd1383	: data1 <= weights[1383];
				12'd1384	: data1 <= weights[1384];
				12'd1385	: data1 <= weights[1385];
				12'd1386	: data1 <= weights[1386];
				12'd1387	: data1 <= weights[1387];
				12'd1388	: data1 <= weights[1388];
				12'd1389	: data1 <= weights[1389];
				12'd1390	: data1 <= weights[1390];
				12'd1391	: data1 <= weights[1391];
				12'd1392	: data1 <= weights[1392];
				12'd1393	: data1 <= weights[1393];
				12'd1394	: data1 <= weights[1394];
				12'd1395	: data1 <= weights[1395];
				12'd1396	: data1 <= weights[1396];
				12'd1397	: data1 <= weights[1397];
				12'd1398	: data1 <= weights[1398];
				12'd1399	: data1 <= weights[1399];
				12'd1400	: data1 <= weights[1400];
				12'd1401	: data1 <= weights[1401];
				12'd1402	: data1 <= weights[1402];
				12'd1403	: data1 <= weights[1403];
				12'd1404	: data1 <= weights[1404];
				12'd1405	: data1 <= weights[1405];
				12'd1406	: data1 <= weights[1406];
				12'd1407	: data1 <= weights[1407];
				12'd1408	: data1 <= weights[1408];
				12'd1409	: data1 <= weights[1409];
				12'd1410	: data1 <= weights[1410];
				12'd1411	: data1 <= weights[1411];
				12'd1412	: data1 <= weights[1412];
				12'd1413	: data1 <= weights[1413];
				12'd1414	: data1 <= weights[1414];
				12'd1415	: data1 <= weights[1415];
				12'd1416	: data1 <= weights[1416];
				12'd1417	: data1 <= weights[1417];
				12'd1418	: data1 <= weights[1418];
				12'd1419	: data1 <= weights[1419];
				12'd1420	: data1 <= weights[1420];
				12'd1421	: data1 <= weights[1421];
				12'd1422	: data1 <= weights[1422];
				12'd1423	: data1 <= weights[1423];
				12'd1424	: data1 <= weights[1424];
				12'd1425	: data1 <= weights[1425];
				12'd1426	: data1 <= weights[1426];
				12'd1427	: data1 <= weights[1427];
				12'd1428	: data1 <= weights[1428];
				12'd1429	: data1 <= weights[1429];
				12'd1430	: data1 <= weights[1430];
				12'd1431	: data1 <= weights[1431];
				12'd1432	: data1 <= weights[1432];
				12'd1433	: data1 <= weights[1433];
				12'd1434	: data1 <= weights[1434];
				12'd1435	: data1 <= weights[1435];
				12'd1436	: data1 <= weights[1436];
				12'd1437	: data1 <= weights[1437];
				12'd1438	: data1 <= weights[1438];
				12'd1439	: data1 <= weights[1439];
				12'd1440	: data1 <= weights[1440];
				12'd1441	: data1 <= weights[1441];
				12'd1442	: data1 <= weights[1442];
				12'd1443	: data1 <= weights[1443];
				12'd1444	: data1 <= weights[1444];
				12'd1445	: data1 <= weights[1445];
				12'd1446	: data1 <= weights[1446];
				12'd1447	: data1 <= weights[1447];
				12'd1448	: data1 <= weights[1448];
				12'd1449	: data1 <= weights[1449];
				12'd1450	: data1 <= weights[1450];
				12'd1451	: data1 <= weights[1451];
				12'd1452	: data1 <= weights[1452];
				12'd1453	: data1 <= weights[1453];
				12'd1454	: data1 <= weights[1454];
				12'd1455	: data1 <= weights[1455];
				12'd1456	: data1 <= weights[1456];
				12'd1457	: data1 <= weights[1457];
				12'd1458	: data1 <= weights[1458];
				12'd1459	: data1 <= weights[1459];
				12'd1460	: data1 <= weights[1460];
				12'd1461	: data1 <= weights[1461];
				12'd1462	: data1 <= weights[1462];
				12'd1463	: data1 <= weights[1463];
				12'd1464	: data1 <= weights[1464];
				12'd1465	: data1 <= weights[1465];
				12'd1466	: data1 <= weights[1466];
				12'd1467	: data1 <= weights[1467];
				12'd1468	: data1 <= weights[1468];
				12'd1469	: data1 <= weights[1469];
				12'd1470	: data1 <= weights[1470];
				12'd1471	: data1 <= weights[1471];
				12'd1472	: data1 <= weights[1472];
				12'd1473	: data1 <= weights[1473];
				12'd1474	: data1 <= weights[1474];
				12'd1475	: data1 <= weights[1475];
				12'd1476	: data1 <= weights[1476];
				12'd1477	: data1 <= weights[1477];
				12'd1478	: data1 <= weights[1478];
				12'd1479	: data1 <= weights[1479];
				12'd1480	: data1 <= weights[1480];
				12'd1481	: data1 <= weights[1481];
				12'd1482	: data1 <= weights[1482];
				12'd1483	: data1 <= weights[1483];
				12'd1484	: data1 <= weights[1484];
				12'd1485	: data1 <= weights[1485];
				12'd1486	: data1 <= weights[1486];
				12'd1487	: data1 <= weights[1487];
				12'd1488	: data1 <= weights[1488];
				12'd1489	: data1 <= weights[1489];
				12'd1490	: data1 <= weights[1490];
				12'd1491	: data1 <= weights[1491];
				12'd1492	: data1 <= weights[1492];
				12'd1493	: data1 <= weights[1493];
				12'd1494	: data1 <= weights[1494];
				12'd1495	: data1 <= weights[1495];
				12'd1496	: data1 <= weights[1496];
				12'd1497	: data1 <= weights[1497];
				12'd1498	: data1 <= weights[1498];
				12'd1499	: data1 <= weights[1499];
				12'd1500	: data1 <= weights[1500];
				12'd1501	: data1 <= weights[1501];
				12'd1502	: data1 <= weights[1502];
				12'd1503	: data1 <= weights[1503];
				12'd1504	: data1 <= weights[1504];
				12'd1505	: data1 <= weights[1505];
				12'd1506	: data1 <= weights[1506];
				12'd1507	: data1 <= weights[1507];
				12'd1508	: data1 <= weights[1508];
				12'd1509	: data1 <= weights[1509];
				12'd1510	: data1 <= weights[1510];
				12'd1511	: data1 <= weights[1511];
				12'd1512	: data1 <= weights[1512];
				12'd1513	: data1 <= weights[1513];
				12'd1514	: data1 <= weights[1514];
				12'd1515	: data1 <= weights[1515];
				12'd1516	: data1 <= weights[1516];
				12'd1517	: data1 <= weights[1517];
				12'd1518	: data1 <= weights[1518];
				12'd1519	: data1 <= weights[1519];
				12'd1520	: data1 <= weights[1520];
				12'd1521	: data1 <= weights[1521];
				12'd1522	: data1 <= weights[1522];
				12'd1523	: data1 <= weights[1523];
				12'd1524	: data1 <= weights[1524];
				12'd1525	: data1 <= weights[1525];
				12'd1526	: data1 <= weights[1526];
				12'd1527	: data1 <= weights[1527];
				12'd1528	: data1 <= weights[1528];
				12'd1529	: data1 <= weights[1529];
				12'd1530	: data1 <= weights[1530];
				12'd1531	: data1 <= weights[1531];
				12'd1532	: data1 <= weights[1532];
				12'd1533	: data1 <= weights[1533];
				12'd1534	: data1 <= weights[1534];
				12'd1535	: data1 <= weights[1535];
				12'd1536	: data1 <= weights[1536];
				12'd1537	: data1 <= weights[1537];
				12'd1538	: data1 <= weights[1538];
				12'd1539	: data1 <= weights[1539];
				12'd1540	: data1 <= weights[1540];
				12'd1541	: data1 <= weights[1541];
				12'd1542	: data1 <= weights[1542];
				12'd1543	: data1 <= weights[1543];
				12'd1544	: data1 <= weights[1544];
				12'd1545	: data1 <= weights[1545];
				12'd1546	: data1 <= weights[1546];
				12'd1547	: data1 <= weights[1547];
				12'd1548	: data1 <= weights[1548];
				12'd1549	: data1 <= weights[1549];
				12'd1550	: data1 <= weights[1550];
				12'd1551	: data1 <= weights[1551];
				12'd1552	: data1 <= weights[1552];
				12'd1553	: data1 <= weights[1553];
				12'd1554	: data1 <= weights[1554];
				12'd1555	: data1 <= weights[1555];
				12'd1556	: data1 <= weights[1556];
				12'd1557	: data1 <= weights[1557];
				12'd1558	: data1 <= weights[1558];
				12'd1559	: data1 <= weights[1559];
				12'd1560	: data1 <= weights[1560];
				12'd1561	: data1 <= weights[1561];
				12'd1562	: data1 <= weights[1562];
				12'd1563	: data1 <= weights[1563];
				12'd1564	: data1 <= weights[1564];
				12'd1565	: data1 <= weights[1565];
				12'd1566	: data1 <= weights[1566];
				12'd1567	: data1 <= weights[1567];
				12'd1568	: data1 <= weights[1568];
				12'd1569	: data1 <= weights[1569];
				12'd1570	: data1 <= weights[1570];
				12'd1571	: data1 <= weights[1571];
				12'd1572	: data1 <= weights[1572];
				12'd1573	: data1 <= weights[1573];
				12'd1574	: data1 <= weights[1574];
				12'd1575	: data1 <= weights[1575];
				12'd1576	: data1 <= weights[1576];
				12'd1577	: data1 <= weights[1577];
				12'd1578	: data1 <= weights[1578];
				12'd1579	: data1 <= weights[1579];
				12'd1580	: data1 <= weights[1580];
				12'd1581	: data1 <= weights[1581];
				12'd1582	: data1 <= weights[1582];
				12'd1583	: data1 <= weights[1583];
				12'd1584	: data1 <= weights[1584];
				12'd1585	: data1 <= weights[1585];
				12'd1586	: data1 <= weights[1586];
				12'd1587	: data1 <= weights[1587];
				12'd1588	: data1 <= weights[1588];
				12'd1589	: data1 <= weights[1589];
				12'd1590	: data1 <= weights[1590];
				12'd1591	: data1 <= weights[1591];
				12'd1592	: data1 <= weights[1592];
				12'd1593	: data1 <= weights[1593];
				12'd1594	: data1 <= weights[1594];
				12'd1595	: data1 <= weights[1595];
				12'd1596	: data1 <= weights[1596];
				12'd1597	: data1 <= weights[1597];
				12'd1598	: data1 <= weights[1598];
				12'd1599	: data1 <= weights[1599];
				12'd1600	: data1 <= weights[1600];
				12'd1601	: data1 <= weights[1601];
				12'd1602	: data1 <= weights[1602];
				12'd1603	: data1 <= weights[1603];
				12'd1604	: data1 <= weights[1604];
				12'd1605	: data1 <= weights[1605];
				12'd1606	: data1 <= weights[1606];
				12'd1607	: data1 <= weights[1607];
				12'd1608	: data1 <= weights[1608];
				12'd1609	: data1 <= weights[1609];
				12'd1610	: data1 <= weights[1610];
				12'd1611	: data1 <= weights[1611];
				12'd1612	: data1 <= weights[1612];
				12'd1613	: data1 <= weights[1613];
				12'd1614	: data1 <= weights[1614];
				12'd1615	: data1 <= weights[1615];
				12'd1616	: data1 <= weights[1616];
				12'd1617	: data1 <= weights[1617];
				12'd1618	: data1 <= weights[1618];
				12'd1619	: data1 <= weights[1619];
				12'd1620	: data1 <= weights[1620];
				12'd1621	: data1 <= weights[1621];
				12'd1622	: data1 <= weights[1622];
				12'd1623	: data1 <= weights[1623];
				12'd1624	: data1 <= weights[1624];
				12'd1625	: data1 <= weights[1625];
				12'd1626	: data1 <= weights[1626];
				12'd1627	: data1 <= weights[1627];
				12'd1628	: data1 <= weights[1628];
				12'd1629	: data1 <= weights[1629];
				12'd1630	: data1 <= weights[1630];
				12'd1631	: data1 <= weights[1631];
				12'd1632	: data1 <= weights[1632];
				12'd1633	: data1 <= weights[1633];
				12'd1634	: data1 <= weights[1634];
				12'd1635	: data1 <= weights[1635];
				12'd1636	: data1 <= weights[1636];
				12'd1637	: data1 <= weights[1637];
				12'd1638	: data1 <= weights[1638];
				12'd1639	: data1 <= weights[1639];
				12'd1640	: data1 <= weights[1640];
				12'd1641	: data1 <= weights[1641];
				12'd1642	: data1 <= weights[1642];
				12'd1643	: data1 <= weights[1643];
				12'd1644	: data1 <= weights[1644];
				12'd1645	: data1 <= weights[1645];
				12'd1646	: data1 <= weights[1646];
				12'd1647	: data1 <= weights[1647];
				12'd1648	: data1 <= weights[1648];
				12'd1649	: data1 <= weights[1649];
				12'd1650	: data1 <= weights[1650];
				12'd1651	: data1 <= weights[1651];
				12'd1652	: data1 <= weights[1652];
				12'd1653	: data1 <= weights[1653];
				12'd1654	: data1 <= weights[1654];
				12'd1655	: data1 <= weights[1655];
				12'd1656	: data1 <= weights[1656];
				12'd1657	: data1 <= weights[1657];
				12'd1658	: data1 <= weights[1658];
				12'd1659	: data1 <= weights[1659];
				12'd1660	: data1 <= weights[1660];
				12'd1661	: data1 <= weights[1661];
				12'd1662	: data1 <= weights[1662];
				12'd1663	: data1 <= weights[1663];
				12'd1664	: data1 <= weights[1664];
				12'd1665	: data1 <= weights[1665];
				12'd1666	: data1 <= weights[1666];
				12'd1667	: data1 <= weights[1667];
				12'd1668	: data1 <= weights[1668];
				12'd1669	: data1 <= weights[1669];
				12'd1670	: data1 <= weights[1670];
				12'd1671	: data1 <= weights[1671];
				12'd1672	: data1 <= weights[1672];
				12'd1673	: data1 <= weights[1673];
				12'd1674	: data1 <= weights[1674];
				12'd1675	: data1 <= weights[1675];
				12'd1676	: data1 <= weights[1676];
				12'd1677	: data1 <= weights[1677];
				12'd1678	: data1 <= weights[1678];
				12'd1679	: data1 <= weights[1679];
				12'd1680	: data1 <= weights[1680];
				12'd1681	: data1 <= weights[1681];
				12'd1682	: data1 <= weights[1682];
				12'd1683	: data1 <= weights[1683];
				12'd1684	: data1 <= weights[1684];
				12'd1685	: data1 <= weights[1685];
				12'd1686	: data1 <= weights[1686];
				12'd1687	: data1 <= weights[1687];
				12'd1688	: data1 <= weights[1688];
				12'd1689	: data1 <= weights[1689];
				12'd1690	: data1 <= weights[1690];
				12'd1691	: data1 <= weights[1691];
				12'd1692	: data1 <= weights[1692];
				12'd1693	: data1 <= weights[1693];
				12'd1694	: data1 <= weights[1694];
				12'd1695	: data1 <= weights[1695];
				12'd1696	: data1 <= weights[1696];
				12'd1697	: data1 <= weights[1697];
				12'd1698	: data1 <= weights[1698];
				12'd1699	: data1 <= weights[1699];
				12'd1700	: data1 <= weights[1700];
				12'd1701	: data1 <= weights[1701];
				12'd1702	: data1 <= weights[1702];
				12'd1703	: data1 <= weights[1703];
				12'd1704	: data1 <= weights[1704];
				12'd1705	: data1 <= weights[1705];
				12'd1706	: data1 <= weights[1706];
				12'd1707	: data1 <= weights[1707];
				12'd1708	: data1 <= weights[1708];
				12'd1709	: data1 <= weights[1709];
				12'd1710	: data1 <= weights[1710];
				12'd1711	: data1 <= weights[1711];
				12'd1712	: data1 <= weights[1712];
				12'd1713	: data1 <= weights[1713];
				12'd1714	: data1 <= weights[1714];
				12'd1715	: data1 <= weights[1715];
				12'd1716	: data1 <= weights[1716];
				12'd1717	: data1 <= weights[1717];
				12'd1718	: data1 <= weights[1718];
				12'd1719	: data1 <= weights[1719];
				12'd1720	: data1 <= weights[1720];
				12'd1721	: data1 <= weights[1721];
				12'd1722	: data1 <= weights[1722];
				12'd1723	: data1 <= weights[1723];
				12'd1724	: data1 <= weights[1724];
				12'd1725	: data1 <= weights[1725];
				12'd1726	: data1 <= weights[1726];
				12'd1727	: data1 <= weights[1727];
				12'd1728	: data1 <= weights[1728];
				12'd1729	: data1 <= weights[1729];
				12'd1730	: data1 <= weights[1730];
				12'd1731	: data1 <= weights[1731];
				12'd1732	: data1 <= weights[1732];
				12'd1733	: data1 <= weights[1733];
				12'd1734	: data1 <= weights[1734];
				12'd1735	: data1 <= weights[1735];
				12'd1736	: data1 <= weights[1736];
				12'd1737	: data1 <= weights[1737];
				12'd1738	: data1 <= weights[1738];
				12'd1739	: data1 <= weights[1739];
				12'd1740	: data1 <= weights[1740];
				12'd1741	: data1 <= weights[1741];
				12'd1742	: data1 <= weights[1742];
				12'd1743	: data1 <= weights[1743];
				12'd1744	: data1 <= weights[1744];
				12'd1745	: data1 <= weights[1745];
				12'd1746	: data1 <= weights[1746];
				12'd1747	: data1 <= weights[1747];
				12'd1748	: data1 <= weights[1748];
				12'd1749	: data1 <= weights[1749];
				12'd1750	: data1 <= weights[1750];
				12'd1751	: data1 <= weights[1751];
				12'd1752	: data1 <= weights[1752];
				12'd1753	: data1 <= weights[1753];
				12'd1754	: data1 <= weights[1754];
				12'd1755	: data1 <= weights[1755];
				12'd1756	: data1 <= weights[1756];
				12'd1757	: data1 <= weights[1757];
				12'd1758	: data1 <= weights[1758];
				12'd1759	: data1 <= weights[1759];
				12'd1760	: data1 <= weights[1760];
				12'd1761	: data1 <= weights[1761];
				12'd1762	: data1 <= weights[1762];
				12'd1763	: data1 <= weights[1763];
				12'd1764	: data1 <= weights[1764];
				12'd1765	: data1 <= weights[1765];
				12'd1766	: data1 <= weights[1766];
				12'd1767	: data1 <= weights[1767];
				12'd1768	: data1 <= weights[1768];
				12'd1769	: data1 <= weights[1769];
				12'd1770	: data1 <= weights[1770];
				12'd1771	: data1 <= weights[1771];
				12'd1772	: data1 <= weights[1772];
				12'd1773	: data1 <= weights[1773];
				12'd1774	: data1 <= weights[1774];
				12'd1775	: data1 <= weights[1775];
				12'd1776	: data1 <= weights[1776];
				12'd1777	: data1 <= weights[1777];
				12'd1778	: data1 <= weights[1778];
				12'd1779	: data1 <= weights[1779];
				12'd1780	: data1 <= weights[1780];
				12'd1781	: data1 <= weights[1781];
				12'd1782	: data1 <= weights[1782];
				12'd1783	: data1 <= weights[1783];
				12'd1784	: data1 <= weights[1784];
				12'd1785	: data1 <= weights[1785];
				12'd1786	: data1 <= weights[1786];
				12'd1787	: data1 <= weights[1787];
				12'd1788	: data1 <= weights[1788];
				12'd1789	: data1 <= weights[1789];
				12'd1790	: data1 <= weights[1790];
				12'd1791	: data1 <= weights[1791];
				12'd1792	: data1 <= weights[1792];
				12'd1793	: data1 <= weights[1793];
				12'd1794	: data1 <= weights[1794];
				12'd1795	: data1 <= weights[1795];
				12'd1796	: data1 <= weights[1796];
				12'd1797	: data1 <= weights[1797];
				12'd1798	: data1 <= weights[1798];
				12'd1799	: data1 <= weights[1799];
				12'd1800	: data1 <= weights[1800];
				12'd1801	: data1 <= weights[1801];
				12'd1802	: data1 <= weights[1802];
				12'd1803	: data1 <= weights[1803];
				12'd1804	: data1 <= weights[1804];
				12'd1805	: data1 <= weights[1805];
				12'd1806	: data1 <= weights[1806];
				12'd1807	: data1 <= weights[1807];
				12'd1808	: data1 <= weights[1808];
				12'd1809	: data1 <= weights[1809];
				12'd1810	: data1 <= weights[1810];
				12'd1811	: data1 <= weights[1811];
				12'd1812	: data1 <= weights[1812];
				12'd1813	: data1 <= weights[1813];
				12'd1814	: data1 <= weights[1814];
				12'd1815	: data1 <= weights[1815];
				12'd1816	: data1 <= weights[1816];
				12'd1817	: data1 <= weights[1817];
				12'd1818	: data1 <= weights[1818];
				12'd1819	: data1 <= weights[1819];
				12'd1820	: data1 <= weights[1820];
				12'd1821	: data1 <= weights[1821];
				12'd1822	: data1 <= weights[1822];
				12'd1823	: data1 <= weights[1823];
				12'd1824	: data1 <= weights[1824];
				12'd1825	: data1 <= weights[1825];
				12'd1826	: data1 <= weights[1826];
				12'd1827	: data1 <= weights[1827];
				12'd1828	: data1 <= weights[1828];
				12'd1829	: data1 <= weights[1829];
				12'd1830	: data1 <= weights[1830];
				12'd1831	: data1 <= weights[1831];
				12'd1832	: data1 <= weights[1832];
				12'd1833	: data1 <= weights[1833];
				12'd1834	: data1 <= weights[1834];
				12'd1835	: data1 <= weights[1835];
				12'd1836	: data1 <= weights[1836];
				12'd1837	: data1 <= weights[1837];
				12'd1838	: data1 <= weights[1838];
				12'd1839	: data1 <= weights[1839];
				12'd1840	: data1 <= weights[1840];
				12'd1841	: data1 <= weights[1841];
				12'd1842	: data1 <= weights[1842];
				12'd1843	: data1 <= weights[1843];
				12'd1844	: data1 <= weights[1844];
				12'd1845	: data1 <= weights[1845];
				12'd1846	: data1 <= weights[1846];
				12'd1847	: data1 <= weights[1847];
				12'd1848	: data1 <= weights[1848];
				12'd1849	: data1 <= weights[1849];
				12'd1850	: data1 <= weights[1850];
				12'd1851	: data1 <= weights[1851];
				12'd1852	: data1 <= weights[1852];
				12'd1853	: data1 <= weights[1853];
				12'd1854	: data1 <= weights[1854];
				12'd1855	: data1 <= weights[1855];
				12'd1856	: data1 <= weights[1856];
				12'd1857	: data1 <= weights[1857];
				12'd1858	: data1 <= weights[1858];
				12'd1859	: data1 <= weights[1859];
				12'd1860	: data1 <= weights[1860];
				12'd1861	: data1 <= weights[1861];
				12'd1862	: data1 <= weights[1862];
				12'd1863	: data1 <= weights[1863];
				12'd1864	: data1 <= weights[1864];
				12'd1865	: data1 <= weights[1865];
				12'd1866	: data1 <= weights[1866];
				12'd1867	: data1 <= weights[1867];
				12'd1868	: data1 <= weights[1868];
				12'd1869	: data1 <= weights[1869];
				12'd1870	: data1 <= weights[1870];
				12'd1871	: data1 <= weights[1871];
				12'd1872	: data1 <= weights[1872];
				12'd1873	: data1 <= weights[1873];
				12'd1874	: data1 <= weights[1874];
				12'd1875	: data1 <= weights[1875];
				12'd1876	: data1 <= weights[1876];
				12'd1877	: data1 <= weights[1877];
				12'd1878	: data1 <= weights[1878];
				12'd1879	: data1 <= weights[1879];
				12'd1880	: data1 <= weights[1880];
				12'd1881	: data1 <= weights[1881];
				12'd1882	: data1 <= weights[1882];
				12'd1883	: data1 <= weights[1883];
				12'd1884	: data1 <= weights[1884];
				12'd1885	: data1 <= weights[1885];
				12'd1886	: data1 <= weights[1886];
				12'd1887	: data1 <= weights[1887];
				12'd1888	: data1 <= weights[1888];
				12'd1889	: data1 <= weights[1889];
				12'd1890	: data1 <= weights[1890];
				12'd1891	: data1 <= weights[1891];
				12'd1892	: data1 <= weights[1892];
				12'd1893	: data1 <= weights[1893];
				12'd1894	: data1 <= weights[1894];
				12'd1895	: data1 <= weights[1895];
				12'd1896	: data1 <= weights[1896];
				12'd1897	: data1 <= weights[1897];
				12'd1898	: data1 <= weights[1898];
				12'd1899	: data1 <= weights[1899];
				12'd1900	: data1 <= weights[1900];
				12'd1901	: data1 <= weights[1901];
				12'd1902	: data1 <= weights[1902];
				12'd1903	: data1 <= weights[1903];
				12'd1904	: data1 <= weights[1904];
				12'd1905	: data1 <= weights[1905];
				12'd1906	: data1 <= weights[1906];
				12'd1907	: data1 <= weights[1907];
				12'd1908	: data1 <= weights[1908];
				12'd1909	: data1 <= weights[1909];
				12'd1910	: data1 <= weights[1910];
				12'd1911	: data1 <= weights[1911];
				12'd1912	: data1 <= weights[1912];
				12'd1913	: data1 <= weights[1913];
				12'd1914	: data1 <= weights[1914];
				12'd1915	: data1 <= weights[1915];
				12'd1916	: data1 <= weights[1916];
				12'd1917	: data1 <= weights[1917];
				12'd1918	: data1 <= weights[1918];
				12'd1919	: data1 <= weights[1919];
				12'd1920	: data1 <= weights[1920];
				12'd1921	: data1 <= weights[1921];
				12'd1922	: data1 <= weights[1922];
				12'd1923	: data1 <= weights[1923];
				12'd1924	: data1 <= weights[1924];
				12'd1925	: data1 <= weights[1925];
				12'd1926	: data1 <= weights[1926];
				12'd1927	: data1 <= weights[1927];
				12'd1928	: data1 <= weights[1928];
				12'd1929	: data1 <= weights[1929];
				12'd1930	: data1 <= weights[1930];
				12'd1931	: data1 <= weights[1931];
				12'd1932	: data1 <= weights[1932];
				12'd1933	: data1 <= weights[1933];
				12'd1934	: data1 <= weights[1934];
				12'd1935	: data1 <= weights[1935];
				12'd1936	: data1 <= weights[1936];
				12'd1937	: data1 <= weights[1937];
				12'd1938	: data1 <= weights[1938];
				12'd1939	: data1 <= weights[1939];
				12'd1940	: data1 <= weights[1940];
				12'd1941	: data1 <= weights[1941];
				12'd1942	: data1 <= weights[1942];
				12'd1943	: data1 <= weights[1943];
				12'd1944	: data1 <= weights[1944];
				12'd1945	: data1 <= weights[1945];
				12'd1946	: data1 <= weights[1946];
				12'd1947	: data1 <= weights[1947];
				12'd1948	: data1 <= weights[1948];
				12'd1949	: data1 <= weights[1949];
				12'd1950	: data1 <= weights[1950];
				12'd1951	: data1 <= weights[1951];
				12'd1952	: data1 <= weights[1952];
				12'd1953	: data1 <= weights[1953];
				12'd1954	: data1 <= weights[1954];
				12'd1955	: data1 <= weights[1955];
				12'd1956	: data1 <= weights[1956];
				12'd1957	: data1 <= weights[1957];
				12'd1958	: data1 <= weights[1958];
				12'd1959	: data1 <= weights[1959];
				12'd1960	: data1 <= weights[1960];
				12'd1961	: data1 <= weights[1961];
				12'd1962	: data1 <= weights[1962];
				12'd1963	: data1 <= weights[1963];
				12'd1964	: data1 <= weights[1964];
				12'd1965	: data1 <= weights[1965];
				12'd1966	: data1 <= weights[1966];
				12'd1967	: data1 <= weights[1967];
				12'd1968	: data1 <= weights[1968];
				12'd1969	: data1 <= weights[1969];
				12'd1970	: data1 <= weights[1970];
				12'd1971	: data1 <= weights[1971];
				12'd1972	: data1 <= weights[1972];
				12'd1973	: data1 <= weights[1973];
				12'd1974	: data1 <= weights[1974];
				12'd1975	: data1 <= weights[1975];
				12'd1976	: data1 <= weights[1976];
				12'd1977	: data1 <= weights[1977];
				12'd1978	: data1 <= weights[1978];
				12'd1979	: data1 <= weights[1979];
				12'd1980	: data1 <= weights[1980];
				12'd1981	: data1 <= weights[1981];
				12'd1982	: data1 <= weights[1982];
				12'd1983	: data1 <= weights[1983];
				12'd1984	: data1 <= weights[1984];
				12'd1985	: data1 <= weights[1985];
				12'd1986	: data1 <= weights[1986];
				12'd1987	: data1 <= weights[1987];
				12'd1988	: data1 <= weights[1988];
				12'd1989	: data1 <= weights[1989];
				12'd1990	: data1 <= weights[1990];
				12'd1991	: data1 <= weights[1991];
				12'd1992	: data1 <= weights[1992];
				12'd1993	: data1 <= weights[1993];
				12'd1994	: data1 <= weights[1994];
				12'd1995	: data1 <= weights[1995];
				12'd1996	: data1 <= weights[1996];
				12'd1997	: data1 <= weights[1997];
				12'd1998	: data1 <= weights[1998];
				12'd1999	: data1 <= weights[1999];
				12'd2000	: data1 <= weights[2000];
				12'd2001	: data1 <= weights[2001];
				12'd2002	: data1 <= weights[2002];
				12'd2003	: data1 <= weights[2003];
				12'd2004	: data1 <= weights[2004];
				12'd2005	: data1 <= weights[2005];
				12'd2006	: data1 <= weights[2006];
				12'd2007	: data1 <= weights[2007];
				12'd2008	: data1 <= weights[2008];
				12'd2009	: data1 <= weights[2009];
				12'd2010	: data1 <= weights[2010];
				12'd2011	: data1 <= weights[2011];
				12'd2012	: data1 <= weights[2012];
				12'd2013	: data1 <= weights[2013];
				12'd2014	: data1 <= weights[2014];
				12'd2015	: data1 <= weights[2015];
				12'd2016	: data1 <= weights[2016];
				12'd2017	: data1 <= weights[2017];
				12'd2018	: data1 <= weights[2018];
				12'd2019	: data1 <= weights[2019];
				12'd2020	: data1 <= weights[2020];
				12'd2021	: data1 <= weights[2021];
				12'd2022	: data1 <= weights[2022];
				12'd2023	: data1 <= weights[2023];
				12'd2024	: data1 <= weights[2024];
				12'd2025	: data1 <= weights[2025];
				12'd2026	: data1 <= weights[2026];
				12'd2027	: data1 <= weights[2027];
				12'd2028	: data1 <= weights[2028];
				12'd2029	: data1 <= weights[2029];
				12'd2030	: data1 <= weights[2030];
				12'd2031	: data1 <= weights[2031];
				12'd2032	: data1 <= weights[2032];
				12'd2033	: data1 <= weights[2033];
				12'd2034	: data1 <= weights[2034];
				12'd2035	: data1 <= weights[2035];
				12'd2036	: data1 <= weights[2036];
				12'd2037	: data1 <= weights[2037];
				12'd2038	: data1 <= weights[2038];
				12'd2039	: data1 <= weights[2039];
				12'd2040	: data1 <= weights[2040];
				12'd2041	: data1 <= weights[2041];
				12'd2042	: data1 <= weights[2042];
				12'd2043	: data1 <= weights[2043];
				12'd2044	: data1 <= weights[2044];
				12'd2045	: data1 <= weights[2045];
				12'd2046	: data1 <= weights[2046];
				12'd2047	: data1 <= weights[2047];
				12'd2048	: data1 <= weights[2048];
				12'd2049	: data1 <= weights[2049];
				12'd2050	: data1 <= weights[2050];
				12'd2051	: data1 <= weights[2051];
				12'd2052	: data1 <= weights[2052];
				12'd2053	: data1 <= weights[2053];
				12'd2054	: data1 <= weights[2054];
				12'd2055	: data1 <= weights[2055];
				12'd2056	: data1 <= weights[2056];
				12'd2057	: data1 <= weights[2057];
				12'd2058	: data1 <= weights[2058];
				12'd2059	: data1 <= weights[2059];
				12'd2060	: data1 <= weights[2060];
				12'd2061	: data1 <= weights[2061];
				12'd2062	: data1 <= weights[2062];
				12'd2063	: data1 <= weights[2063];
				12'd2064	: data1 <= weights[2064];
				12'd2065	: data1 <= weights[2065];
				12'd2066	: data1 <= weights[2066];
				12'd2067	: data1 <= weights[2067];
				12'd2068	: data1 <= weights[2068];
				12'd2069	: data1 <= weights[2069];
				12'd2070	: data1 <= weights[2070];
				12'd2071	: data1 <= weights[2071];
				12'd2072	: data1 <= weights[2072];
				12'd2073	: data1 <= weights[2073];
				12'd2074	: data1 <= weights[2074];
				12'd2075	: data1 <= weights[2075];
				12'd2076	: data1 <= weights[2076];
				12'd2077	: data1 <= weights[2077];
				12'd2078	: data1 <= weights[2078];
				12'd2079	: data1 <= weights[2079];
				12'd2080	: data1 <= weights[2080];
				12'd2081	: data1 <= weights[2081];
				12'd2082	: data1 <= weights[2082];
				12'd2083	: data1 <= weights[2083];
				12'd2084	: data1 <= weights[2084];
				12'd2085	: data1 <= weights[2085];
				12'd2086	: data1 <= weights[2086];
				12'd2087	: data1 <= weights[2087];
				12'd2088	: data1 <= weights[2088];
				12'd2089	: data1 <= weights[2089];
				12'd2090	: data1 <= weights[2090];
				12'd2091	: data1 <= weights[2091];
				12'd2092	: data1 <= weights[2092];
				12'd2093	: data1 <= weights[2093];
				12'd2094	: data1 <= weights[2094];
				12'd2095	: data1 <= weights[2095];
				12'd2096	: data1 <= weights[2096];
				12'd2097	: data1 <= weights[2097];
				12'd2098	: data1 <= weights[2098];
				12'd2099	: data1 <= weights[2099];
				12'd2100	: data1 <= weights[2100];
				12'd2101	: data1 <= weights[2101];
				12'd2102	: data1 <= weights[2102];
				12'd2103	: data1 <= weights[2103];
				12'd2104	: data1 <= weights[2104];
				12'd2105	: data1 <= weights[2105];
				12'd2106	: data1 <= weights[2106];
				12'd2107	: data1 <= weights[2107];
				12'd2108	: data1 <= weights[2108];
				12'd2109	: data1 <= weights[2109];
				12'd2110	: data1 <= weights[2110];
				12'd2111	: data1 <= weights[2111];
				12'd2112	: data1 <= weights[2112];
				12'd2113	: data1 <= weights[2113];
				12'd2114	: data1 <= weights[2114];
				12'd2115	: data1 <= weights[2115];
				12'd2116	: data1 <= weights[2116];
				12'd2117	: data1 <= weights[2117];
				12'd2118	: data1 <= weights[2118];
				12'd2119	: data1 <= weights[2119];
				12'd2120	: data1 <= weights[2120];
				12'd2121	: data1 <= weights[2121];
				12'd2122	: data1 <= weights[2122];
				12'd2123	: data1 <= weights[2123];
				12'd2124	: data1 <= weights[2124];
				12'd2125	: data1 <= weights[2125];
				12'd2126	: data1 <= weights[2126];
				12'd2127	: data1 <= weights[2127];
				12'd2128	: data1 <= weights[2128];
				12'd2129	: data1 <= weights[2129];
				12'd2130	: data1 <= weights[2130];
				12'd2131	: data1 <= weights[2131];
				12'd2132	: data1 <= weights[2132];
				12'd2133	: data1 <= weights[2133];
				12'd2134	: data1 <= weights[2134];
				12'd2135	: data1 <= weights[2135];
				12'd2136	: data1 <= weights[2136];
				12'd2137	: data1 <= weights[2137];
				12'd2138	: data1 <= weights[2138];
				12'd2139	: data1 <= weights[2139];
				12'd2140	: data1 <= weights[2140];
				12'd2141	: data1 <= weights[2141];
				12'd2142	: data1 <= weights[2142];
				12'd2143	: data1 <= weights[2143];
				12'd2144	: data1 <= weights[2144];
				12'd2145	: data1 <= weights[2145];
				12'd2146	: data1 <= weights[2146];
				12'd2147	: data1 <= weights[2147];
				12'd2148	: data1 <= weights[2148];
				12'd2149	: data1 <= weights[2149];
				12'd2150	: data1 <= weights[2150];
				12'd2151	: data1 <= weights[2151];
				12'd2152	: data1 <= weights[2152];
				12'd2153	: data1 <= weights[2153];
				12'd2154	: data1 <= weights[2154];
				12'd2155	: data1 <= weights[2155];
				12'd2156	: data1 <= weights[2156];
				12'd2157	: data1 <= weights[2157];
				12'd2158	: data1 <= weights[2158];
				12'd2159	: data1 <= weights[2159];
				12'd2160	: data1 <= weights[2160];
				12'd2161	: data1 <= weights[2161];
				12'd2162	: data1 <= weights[2162];
				12'd2163	: data1 <= weights[2163];
				12'd2164	: data1 <= weights[2164];
				12'd2165	: data1 <= weights[2165];
				12'd2166	: data1 <= weights[2166];
				12'd2167	: data1 <= weights[2167];
				12'd2168	: data1 <= weights[2168];
				12'd2169	: data1 <= weights[2169];
				12'd2170	: data1 <= weights[2170];
				12'd2171	: data1 <= weights[2171];
				12'd2172	: data1 <= weights[2172];
				12'd2173	: data1 <= weights[2173];
				12'd2174	: data1 <= weights[2174];
				12'd2175	: data1 <= weights[2175];
				12'd2176	: data1 <= weights[2176];
				12'd2177	: data1 <= weights[2177];
				12'd2178	: data1 <= weights[2178];
				12'd2179	: data1 <= weights[2179];
				12'd2180	: data1 <= weights[2180];
				12'd2181	: data1 <= weights[2181];
				12'd2182	: data1 <= weights[2182];
				12'd2183	: data1 <= weights[2183];
				12'd2184	: data1 <= weights[2184];
				12'd2185	: data1 <= weights[2185];
				12'd2186	: data1 <= weights[2186];
				12'd2187	: data1 <= weights[2187];
				12'd2188	: data1 <= weights[2188];
				12'd2189	: data1 <= weights[2189];
				12'd2190	: data1 <= weights[2190];
				12'd2191	: data1 <= weights[2191];
				12'd2192	: data1 <= weights[2192];
				12'd2193	: data1 <= weights[2193];
				12'd2194	: data1 <= weights[2194];
				12'd2195	: data1 <= weights[2195];
				12'd2196	: data1 <= weights[2196];
				12'd2197	: data1 <= weights[2197];
				12'd2198	: data1 <= weights[2198];
				12'd2199	: data1 <= weights[2199];
				12'd2200	: data1 <= weights[2200];
				12'd2201	: data1 <= weights[2201];
				12'd2202	: data1 <= weights[2202];
				12'd2203	: data1 <= weights[2203];
				12'd2204	: data1 <= weights[2204];
				12'd2205	: data1 <= weights[2205];
				12'd2206	: data1 <= weights[2206];
				12'd2207	: data1 <= weights[2207];
				12'd2208	: data1 <= weights[2208];
				12'd2209	: data1 <= weights[2209];
				12'd2210	: data1 <= weights[2210];
				12'd2211	: data1 <= weights[2211];
				12'd2212	: data1 <= weights[2212];
				12'd2213	: data1 <= weights[2213];
				12'd2214	: data1 <= weights[2214];
				12'd2215	: data1 <= weights[2215];
				12'd2216	: data1 <= weights[2216];
				12'd2217	: data1 <= weights[2217];
				12'd2218	: data1 <= weights[2218];
				12'd2219	: data1 <= weights[2219];
				12'd2220	: data1 <= weights[2220];
				12'd2221	: data1 <= weights[2221];
				12'd2222	: data1 <= weights[2222];
				12'd2223	: data1 <= weights[2223];
				12'd2224	: data1 <= weights[2224];
				12'd2225	: data1 <= weights[2225];
				12'd2226	: data1 <= weights[2226];
				12'd2227	: data1 <= weights[2227];
				12'd2228	: data1 <= weights[2228];
				12'd2229	: data1 <= weights[2229];
				12'd2230	: data1 <= weights[2230];
				12'd2231	: data1 <= weights[2231];
				12'd2232	: data1 <= weights[2232];
				12'd2233	: data1 <= weights[2233];
				12'd2234	: data1 <= weights[2234];
				12'd2235	: data1 <= weights[2235];
				12'd2236	: data1 <= weights[2236];
				12'd2237	: data1 <= weights[2237];
				12'd2238	: data1 <= weights[2238];
				12'd2239	: data1 <= weights[2239];
				12'd2240	: data1 <= weights[2240];
				12'd2241	: data1 <= weights[2241];
				12'd2242	: data1 <= weights[2242];
				12'd2243	: data1 <= weights[2243];
				12'd2244	: data1 <= weights[2244];
				12'd2245	: data1 <= weights[2245];
				12'd2246	: data1 <= weights[2246];
				12'd2247	: data1 <= weights[2247];
				12'd2248	: data1 <= weights[2248];
				12'd2249	: data1 <= weights[2249];
				12'd2250	: data1 <= weights[2250];
				12'd2251	: data1 <= weights[2251];
				12'd2252	: data1 <= weights[2252];
				12'd2253	: data1 <= weights[2253];
				12'd2254	: data1 <= weights[2254];
				12'd2255	: data1 <= weights[2255];
				12'd2256	: data1 <= weights[2256];
				12'd2257	: data1 <= weights[2257];
				12'd2258	: data1 <= weights[2258];
				12'd2259	: data1 <= weights[2259];
				12'd2260	: data1 <= weights[2260];
				12'd2261	: data1 <= weights[2261];
				12'd2262	: data1 <= weights[2262];
				12'd2263	: data1 <= weights[2263];
				12'd2264	: data1 <= weights[2264];
				12'd2265	: data1 <= weights[2265];
				12'd2266	: data1 <= weights[2266];
				12'd2267	: data1 <= weights[2267];
				12'd2268	: data1 <= weights[2268];
				12'd2269	: data1 <= weights[2269];
				12'd2270	: data1 <= weights[2270];
				12'd2271	: data1 <= weights[2271];
				12'd2272	: data1 <= weights[2272];
				12'd2273	: data1 <= weights[2273];
				12'd2274	: data1 <= weights[2274];
				12'd2275	: data1 <= weights[2275];
				12'd2276	: data1 <= weights[2276];
				12'd2277	: data1 <= weights[2277];
				12'd2278	: data1 <= weights[2278];
				12'd2279	: data1 <= weights[2279];
				12'd2280	: data1 <= weights[2280];
				12'd2281	: data1 <= weights[2281];
				12'd2282	: data1 <= weights[2282];
				12'd2283	: data1 <= weights[2283];
				12'd2284	: data1 <= weights[2284];
				12'd2285	: data1 <= weights[2285];
				12'd2286	: data1 <= weights[2286];
				12'd2287	: data1 <= weights[2287];
				12'd2288	: data1 <= weights[2288];
				12'd2289	: data1 <= weights[2289];
				12'd2290	: data1 <= weights[2290];
				12'd2291	: data1 <= weights[2291];
				12'd2292	: data1 <= weights[2292];
				12'd2293	: data1 <= weights[2293];
				12'd2294	: data1 <= weights[2294];
				12'd2295	: data1 <= weights[2295];
				12'd2296	: data1 <= weights[2296];
				12'd2297	: data1 <= weights[2297];
				12'd2298	: data1 <= weights[2298];
				12'd2299	: data1 <= weights[2299];
				12'd2300	: data1 <= weights[2300];
				12'd2301	: data1 <= weights[2301];
				12'd2302	: data1 <= weights[2302];
				12'd2303	: data1 <= weights[2303];
				12'd2304	: data1 <= weights[2304];
				12'd2305	: data1 <= weights[2305];
				12'd2306	: data1 <= weights[2306];
				12'd2307	: data1 <= weights[2307];
				12'd2308	: data1 <= weights[2308];
				12'd2309	: data1 <= weights[2309];
				12'd2310	: data1 <= weights[2310];
				12'd2311	: data1 <= weights[2311];
				12'd2312	: data1 <= weights[2312];
				12'd2313	: data1 <= weights[2313];
				12'd2314	: data1 <= weights[2314];
				12'd2315	: data1 <= weights[2315];
				12'd2316	: data1 <= weights[2316];
				12'd2317	: data1 <= weights[2317];
				12'd2318	: data1 <= weights[2318];
				12'd2319	: data1 <= weights[2319];
				12'd2320	: data1 <= weights[2320];
				12'd2321	: data1 <= weights[2321];
				12'd2322	: data1 <= weights[2322];
				12'd2323	: data1 <= weights[2323];
				12'd2324	: data1 <= weights[2324];
				12'd2325	: data1 <= weights[2325];
				12'd2326	: data1 <= weights[2326];
				12'd2327	: data1 <= weights[2327];
				12'd2328	: data1 <= weights[2328];
				12'd2329	: data1 <= weights[2329];
				12'd2330	: data1 <= weights[2330];
				12'd2331	: data1 <= weights[2331];
				12'd2332	: data1 <= weights[2332];
				12'd2333	: data1 <= weights[2333];
				12'd2334	: data1 <= weights[2334];
				12'd2335	: data1 <= weights[2335];
				12'd2336	: data1 <= weights[2336];
				12'd2337	: data1 <= weights[2337];
				12'd2338	: data1 <= weights[2338];
				12'd2339	: data1 <= weights[2339];
				12'd2340	: data1 <= weights[2340];
				12'd2341	: data1 <= weights[2341];
				12'd2342	: data1 <= weights[2342];
				12'd2343	: data1 <= weights[2343];
				12'd2344	: data1 <= weights[2344];
				12'd2345	: data1 <= weights[2345];
				12'd2346	: data1 <= weights[2346];
				12'd2347	: data1 <= weights[2347];
				12'd2348	: data1 <= weights[2348];
				12'd2349	: data1 <= weights[2349];
				12'd2350	: data1 <= weights[2350];
				12'd2351	: data1 <= weights[2351];
				12'd2352	: data1 <= weights[2352];
				12'd2353	: data1 <= weights[2353];
				12'd2354	: data1 <= weights[2354];
				12'd2355	: data1 <= weights[2355];
				12'd2356	: data1 <= weights[2356];
				12'd2357	: data1 <= weights[2357];
				12'd2358	: data1 <= weights[2358];
				12'd2359	: data1 <= weights[2359];
				12'd2360	: data1 <= weights[2360];
				12'd2361	: data1 <= weights[2361];
				12'd2362	: data1 <= weights[2362];
				12'd2363	: data1 <= weights[2363];
				12'd2364	: data1 <= weights[2364];
				12'd2365	: data1 <= weights[2365];
				12'd2366	: data1 <= weights[2366];
				12'd2367	: data1 <= weights[2367];
				12'd2368	: data1 <= weights[2368];
				12'd2369	: data1 <= weights[2369];
				12'd2370	: data1 <= weights[2370];
				12'd2371	: data1 <= weights[2371];
				12'd2372	: data1 <= weights[2372];
				12'd2373	: data1 <= weights[2373];
				12'd2374	: data1 <= weights[2374];
				12'd2375	: data1 <= weights[2375];
				12'd2376	: data1 <= weights[2376];
				12'd2377	: data1 <= weights[2377];
				12'd2378	: data1 <= weights[2378];
				12'd2379	: data1 <= weights[2379];
				12'd2380	: data1 <= weights[2380];
				12'd2381	: data1 <= weights[2381];
				12'd2382	: data1 <= weights[2382];
				12'd2383	: data1 <= weights[2383];
				12'd2384	: data1 <= weights[2384];
				12'd2385	: data1 <= weights[2385];
				12'd2386	: data1 <= weights[2386];
				12'd2387	: data1 <= weights[2387];
				12'd2388	: data1 <= weights[2388];
				12'd2389	: data1 <= weights[2389];
				12'd2390	: data1 <= weights[2390];
				12'd2391	: data1 <= weights[2391];
				12'd2392	: data1 <= weights[2392];
				12'd2393	: data1 <= weights[2393];
				12'd2394	: data1 <= weights[2394];
				12'd2395	: data1 <= weights[2395];
				12'd2396	: data1 <= weights[2396];
				12'd2397	: data1 <= weights[2397];
				12'd2398	: data1 <= weights[2398];
				12'd2399	: data1 <= weights[2399];
				12'd2400	: data1 <= weights[2400];
				12'd2401	: data1 <= weights[2401];
				12'd2402	: data1 <= weights[2402];
				12'd2403	: data1 <= weights[2403];
				12'd2404	: data1 <= weights[2404];
				12'd2405	: data1 <= weights[2405];
				12'd2406	: data1 <= weights[2406];
				12'd2407	: data1 <= weights[2407];
				12'd2408	: data1 <= weights[2408];
				12'd2409	: data1 <= weights[2409];
				12'd2410	: data1 <= weights[2410];
				12'd2411	: data1 <= weights[2411];
				12'd2412	: data1 <= weights[2412];
				12'd2413	: data1 <= weights[2413];
				12'd2414	: data1 <= weights[2414];
				12'd2415	: data1 <= weights[2415];
				12'd2416	: data1 <= weights[2416];
				12'd2417	: data1 <= weights[2417];
				12'd2418	: data1 <= weights[2418];
				12'd2419	: data1 <= weights[2419];
				12'd2420	: data1 <= weights[2420];
				12'd2421	: data1 <= weights[2421];
				12'd2422	: data1 <= weights[2422];
				12'd2423	: data1 <= weights[2423];
				12'd2424	: data1 <= weights[2424];
				12'd2425	: data1 <= weights[2425];
				12'd2426	: data1 <= weights[2426];
				12'd2427	: data1 <= weights[2427];
				12'd2428	: data1 <= weights[2428];
				12'd2429	: data1 <= weights[2429];
				12'd2430	: data1 <= weights[2430];
				12'd2431	: data1 <= weights[2431];
				12'd2432	: data1 <= weights[2432];
				12'd2433	: data1 <= weights[2433];
				12'd2434	: data1 <= weights[2434];
				12'd2435	: data1 <= weights[2435];
				12'd2436	: data1 <= weights[2436];
				12'd2437	: data1 <= weights[2437];
				12'd2438	: data1 <= weights[2438];
				12'd2439	: data1 <= weights[2439];
				12'd2440	: data1 <= weights[2440];
				12'd2441	: data1 <= weights[2441];
				12'd2442	: data1 <= weights[2442];
				12'd2443	: data1 <= weights[2443];
				12'd2444	: data1 <= weights[2444];
				12'd2445	: data1 <= weights[2445];
				12'd2446	: data1 <= weights[2446];
				12'd2447	: data1 <= weights[2447];
				12'd2448	: data1 <= weights[2448];
				12'd2449	: data1 <= weights[2449];
				12'd2450	: data1 <= weights[2450];
				12'd2451	: data1 <= weights[2451];
				12'd2452	: data1 <= weights[2452];
				12'd2453	: data1 <= weights[2453];
				12'd2454	: data1 <= weights[2454];
				12'd2455	: data1 <= weights[2455];
				12'd2456	: data1 <= weights[2456];
				12'd2457	: data1 <= weights[2457];
				12'd2458	: data1 <= weights[2458];
				12'd2459	: data1 <= weights[2459];
				12'd2460	: data1 <= weights[2460];
				12'd2461	: data1 <= weights[2461];
				12'd2462	: data1 <= weights[2462];
				12'd2463	: data1 <= weights[2463];
				12'd2464	: data1 <= weights[2464];
				12'd2465	: data1 <= weights[2465];
				12'd2466	: data1 <= weights[2466];
				12'd2467	: data1 <= weights[2467];
				12'd2468	: data1 <= weights[2468];
				12'd2469	: data1 <= weights[2469];
				12'd2470	: data1 <= weights[2470];
				12'd2471	: data1 <= weights[2471];
				12'd2472	: data1 <= weights[2472];
				12'd2473	: data1 <= weights[2473];
				12'd2474	: data1 <= weights[2474];
				12'd2475	: data1 <= weights[2475];
				12'd2476	: data1 <= weights[2476];
				12'd2477	: data1 <= weights[2477];
				12'd2478	: data1 <= weights[2478];
				12'd2479	: data1 <= weights[2479];
				12'd2480	: data1 <= weights[2480];
				12'd2481	: data1 <= weights[2481];
				12'd2482	: data1 <= weights[2482];
				12'd2483	: data1 <= weights[2483];
				12'd2484	: data1 <= weights[2484];
				12'd2485	: data1 <= weights[2485];
				12'd2486	: data1 <= weights[2486];
				12'd2487	: data1 <= weights[2487];
				12'd2488	: data1 <= weights[2488];
				12'd2489	: data1 <= weights[2489];
				12'd2490	: data1 <= weights[2490];
				12'd2491	: data1 <= weights[2491];
				12'd2492	: data1 <= weights[2492];
				12'd2493	: data1 <= weights[2493];
				12'd2494	: data1 <= weights[2494];
				12'd2495	: data1 <= weights[2495];
				12'd2496	: data1 <= weights[2496];
				12'd2497	: data1 <= weights[2497];
				12'd2498	: data1 <= weights[2498];
				12'd2499	: data1 <= weights[2499];
				12'd2500	: data1 <= weights[2500];
				12'd2501	: data1 <= weights[2501];
				12'd2502	: data1 <= weights[2502];
				12'd2503	: data1 <= weights[2503];
				12'd2504	: data1 <= weights[2504];
				12'd2505	: data1 <= weights[2505];
				12'd2506	: data1 <= weights[2506];
				12'd2507	: data1 <= weights[2507];
				12'd2508	: data1 <= weights[2508];
				12'd2509	: data1 <= weights[2509];
				12'd2510	: data1 <= weights[2510];
				12'd2511	: data1 <= weights[2511];
				12'd2512	: data1 <= weights[2512];
				12'd2513	: data1 <= weights[2513];
				12'd2514	: data1 <= weights[2514];
				12'd2515	: data1 <= weights[2515];
				12'd2516	: data1 <= weights[2516];
				12'd2517	: data1 <= weights[2517];
				12'd2518	: data1 <= weights[2518];
				12'd2519	: data1 <= weights[2519];
				12'd2520	: data1 <= weights[2520];
				12'd2521	: data1 <= weights[2521];
				12'd2522	: data1 <= weights[2522];
				12'd2523	: data1 <= weights[2523];
				12'd2524	: data1 <= weights[2524];
				12'd2525	: data1 <= weights[2525];
				12'd2526	: data1 <= weights[2526];
				12'd2527	: data1 <= weights[2527];
				12'd2528	: data1 <= weights[2528];
				12'd2529	: data1 <= weights[2529];
				12'd2530	: data1 <= weights[2530];
				12'd2531	: data1 <= weights[2531];
				12'd2532	: data1 <= weights[2532];
				12'd2533	: data1 <= weights[2533];
				12'd2534	: data1 <= weights[2534];
				12'd2535	: data1 <= weights[2535];
				12'd2536	: data1 <= weights[2536];
				12'd2537	: data1 <= weights[2537];
				12'd2538	: data1 <= weights[2538];
				12'd2539	: data1 <= weights[2539];
				12'd2540	: data1 <= weights[2540];
				12'd2541	: data1 <= weights[2541];
				12'd2542	: data1 <= weights[2542];
				12'd2543	: data1 <= weights[2543];
				12'd2544	: data1 <= weights[2544];
				12'd2545	: data1 <= weights[2545];
				12'd2546	: data1 <= weights[2546];
				12'd2547	: data1 <= weights[2547];
				12'd2548	: data1 <= weights[2548];
				12'd2549	: data1 <= weights[2549];
				12'd2550	: data1 <= weights[2550];
				12'd2551	: data1 <= weights[2551];
				12'd2552	: data1 <= weights[2552];
				12'd2553	: data1 <= weights[2553];
				12'd2554	: data1 <= weights[2554];
				12'd2555	: data1 <= weights[2555];
				12'd2556	: data1 <= weights[2556];
				12'd2557	: data1 <= weights[2557];
				12'd2558	: data1 <= weights[2558];
				12'd2559	: data1 <= weights[2559];
				12'd2560	: data1 <= weights[2560];
				12'd2561	: data1 <= weights[2561];
				12'd2562	: data1 <= weights[2562];
				12'd2563	: data1 <= weights[2563];
				12'd2564	: data1 <= weights[2564];
				12'd2565	: data1 <= weights[2565];
				12'd2566	: data1 <= weights[2566];
				12'd2567	: data1 <= weights[2567];
				12'd2568	: data1 <= weights[2568];
				12'd2569	: data1 <= weights[2569];
				12'd2570	: data1 <= weights[2570];
				12'd2571	: data1 <= weights[2571];
				12'd2572	: data1 <= weights[2572];
				12'd2573	: data1 <= weights[2573];
				12'd2574	: data1 <= weights[2574];
				12'd2575	: data1 <= weights[2575];
				12'd2576	: data1 <= weights[2576];
				12'd2577	: data1 <= weights[2577];
				12'd2578	: data1 <= weights[2578];
				12'd2579	: data1 <= weights[2579];
				12'd2580	: data1 <= weights[2580];
				12'd2581	: data1 <= weights[2581];
				12'd2582	: data1 <= weights[2582];
				12'd2583	: data1 <= weights[2583];
				12'd2584	: data1 <= weights[2584];
				12'd2585	: data1 <= weights[2585];
				12'd2586	: data1 <= weights[2586];
				12'd2587	: data1 <= weights[2587];
				12'd2588	: data1 <= weights[2588];
				12'd2589	: data1 <= weights[2589];
				12'd2590	: data1 <= weights[2590];
				12'd2591	: data1 <= weights[2591];
				12'd2592	: data1 <= weights[2592];
				12'd2593	: data1 <= weights[2593];
				12'd2594	: data1 <= weights[2594];
				12'd2595	: data1 <= weights[2595];
				12'd2596	: data1 <= weights[2596];
				12'd2597	: data1 <= weights[2597];
				12'd2598	: data1 <= weights[2598];
				12'd2599	: data1 <= weights[2599];
				12'd2600	: data1 <= weights[2600];
				12'd2601	: data1 <= weights[2601];
				12'd2602	: data1 <= weights[2602];
				12'd2603	: data1 <= weights[2603];
				12'd2604	: data1 <= weights[2604];
				12'd2605	: data1 <= weights[2605];
				12'd2606	: data1 <= weights[2606];
				12'd2607	: data1 <= weights[2607];
				12'd2608	: data1 <= weights[2608];
				12'd2609	: data1 <= weights[2609];
				12'd2610	: data1 <= weights[2610];
				12'd2611	: data1 <= weights[2611];
				12'd2612	: data1 <= weights[2612];
				12'd2613	: data1 <= weights[2613];
				12'd2614	: data1 <= weights[2614];
				12'd2615	: data1 <= weights[2615];
				12'd2616	: data1 <= weights[2616];
				12'd2617	: data1 <= weights[2617];
				12'd2618	: data1 <= weights[2618];
				12'd2619	: data1 <= weights[2619];
				12'd2620	: data1 <= weights[2620];
				12'd2621	: data1 <= weights[2621];
				12'd2622	: data1 <= weights[2622];
				12'd2623	: data1 <= weights[2623];
				12'd2624	: data1 <= weights[2624];
				12'd2625	: data1 <= weights[2625];
				12'd2626	: data1 <= weights[2626];
				12'd2627	: data1 <= weights[2627];
				12'd2628	: data1 <= weights[2628];
				12'd2629	: data1 <= weights[2629];
				12'd2630	: data1 <= weights[2630];
				12'd2631	: data1 <= weights[2631];
				12'd2632	: data1 <= weights[2632];
				12'd2633	: data1 <= weights[2633];
				12'd2634	: data1 <= weights[2634];
				12'd2635	: data1 <= weights[2635];
				12'd2636	: data1 <= weights[2636];
				12'd2637	: data1 <= weights[2637];
				12'd2638	: data1 <= weights[2638];
				12'd2639	: data1 <= weights[2639];
				12'd2640	: data1 <= weights[2640];
				12'd2641	: data1 <= weights[2641];
				12'd2642	: data1 <= weights[2642];
				12'd2643	: data1 <= weights[2643];
				12'd2644	: data1 <= weights[2644];
				12'd2645	: data1 <= weights[2645];
				12'd2646	: data1 <= weights[2646];
				12'd2647	: data1 <= weights[2647];
				12'd2648	: data1 <= weights[2648];
				12'd2649	: data1 <= weights[2649];
				12'd2650	: data1 <= weights[2650];
				12'd2651	: data1 <= weights[2651];
				12'd2652	: data1 <= weights[2652];
				12'd2653	: data1 <= weights[2653];
				12'd2654	: data1 <= weights[2654];
				12'd2655	: data1 <= weights[2655];
				12'd2656	: data1 <= weights[2656];
				12'd2657	: data1 <= weights[2657];
				12'd2658	: data1 <= weights[2658];
				12'd2659	: data1 <= weights[2659];
				12'd2660	: data1 <= weights[2660];
				12'd2661	: data1 <= weights[2661];
				12'd2662	: data1 <= weights[2662];
				12'd2663	: data1 <= weights[2663];
				12'd2664	: data1 <= weights[2664];
				12'd2665	: data1 <= weights[2665];
				12'd2666	: data1 <= weights[2666];
				12'd2667	: data1 <= weights[2667];
				12'd2668	: data1 <= weights[2668];
				12'd2669	: data1 <= weights[2669];
				12'd2670	: data1 <= weights[2670];
				12'd2671	: data1 <= weights[2671];
				12'd2672	: data1 <= weights[2672];
				12'd2673	: data1 <= weights[2673];
				12'd2674	: data1 <= weights[2674];
				12'd2675	: data1 <= weights[2675];
				12'd2676	: data1 <= weights[2676];
				12'd2677	: data1 <= weights[2677];
				12'd2678	: data1 <= weights[2678];
				12'd2679	: data1 <= weights[2679];
				12'd2680	: data1 <= weights[2680];
				12'd2681	: data1 <= weights[2681];
				12'd2682	: data1 <= weights[2682];
				12'd2683	: data1 <= weights[2683];
				12'd2684	: data1 <= weights[2684];
				12'd2685	: data1 <= weights[2685];
				12'd2686	: data1 <= weights[2686];
				12'd2687	: data1 <= weights[2687];
				12'd2688	: data1 <= weights[2688];
				12'd2689	: data1 <= weights[2689];
				12'd2690	: data1 <= weights[2690];
				12'd2691	: data1 <= weights[2691];
				12'd2692	: data1 <= weights[2692];
				12'd2693	: data1 <= weights[2693];
				12'd2694	: data1 <= weights[2694];
				12'd2695	: data1 <= weights[2695];
				12'd2696	: data1 <= weights[2696];
				12'd2697	: data1 <= weights[2697];
				12'd2698	: data1 <= weights[2698];
				12'd2699	: data1 <= weights[2699];
				12'd2700	: data1 <= weights[2700];
				12'd2701	: data1 <= weights[2701];
				12'd2702	: data1 <= weights[2702];
				12'd2703	: data1 <= weights[2703];
				12'd2704	: data1 <= weights[2704];
				12'd2705	: data1 <= weights[2705];
				12'd2706	: data1 <= weights[2706];
				12'd2707	: data1 <= weights[2707];
				12'd2708	: data1 <= weights[2708];
				12'd2709	: data1 <= weights[2709];
				12'd2710	: data1 <= weights[2710];
				12'd2711	: data1 <= weights[2711];
				12'd2712	: data1 <= weights[2712];
				12'd2713	: data1 <= weights[2713];
				12'd2714	: data1 <= weights[2714];
				12'd2715	: data1 <= weights[2715];
				12'd2716	: data1 <= weights[2716];
				12'd2717	: data1 <= weights[2717];
				12'd2718	: data1 <= weights[2718];
				12'd2719	: data1 <= weights[2719];
				12'd2720	: data1 <= weights[2720];
				12'd2721	: data1 <= weights[2721];
				12'd2722	: data1 <= weights[2722];
				12'd2723	: data1 <= weights[2723];
				12'd2724	: data1 <= weights[2724];
				12'd2725	: data1 <= weights[2725];
				12'd2726	: data1 <= weights[2726];
				12'd2727	: data1 <= weights[2727];
				12'd2728	: data1 <= weights[2728];
				12'd2729	: data1 <= weights[2729];
				12'd2730	: data1 <= weights[2730];
				12'd2731	: data1 <= weights[2731];
				12'd2732	: data1 <= weights[2732];
				12'd2733	: data1 <= weights[2733];
				12'd2734	: data1 <= weights[2734];
				12'd2735	: data1 <= weights[2735];
				12'd2736	: data1 <= weights[2736];
				12'd2737	: data1 <= weights[2737];
				12'd2738	: data1 <= weights[2738];
				12'd2739	: data1 <= weights[2739];
				12'd2740	: data1 <= weights[2740];
				12'd2741	: data1 <= weights[2741];
				12'd2742	: data1 <= weights[2742];
				12'd2743	: data1 <= weights[2743];
				12'd2744	: data1 <= weights[2744];
				12'd2745	: data1 <= weights[2745];
				12'd2746	: data1 <= weights[2746];
				12'd2747	: data1 <= weights[2747];
				12'd2748	: data1 <= weights[2748];
				12'd2749	: data1 <= weights[2749];
				12'd2750	: data1 <= weights[2750];
				12'd2751	: data1 <= weights[2751];
				12'd2752	: data1 <= weights[2752];
				12'd2753	: data1 <= weights[2753];
				12'd2754	: data1 <= weights[2754];
				12'd2755	: data1 <= weights[2755];
				12'd2756	: data1 <= weights[2756];
				12'd2757	: data1 <= weights[2757];
				12'd2758	: data1 <= weights[2758];
				12'd2759	: data1 <= weights[2759];
				12'd2760	: data1 <= weights[2760];
				12'd2761	: data1 <= weights[2761];
				12'd2762	: data1 <= weights[2762];
				12'd2763	: data1 <= weights[2763];
				12'd2764	: data1 <= weights[2764];
				12'd2765	: data1 <= weights[2765];
				12'd2766	: data1 <= weights[2766];
				12'd2767	: data1 <= weights[2767];
				12'd2768	: data1 <= weights[2768];
				12'd2769	: data1 <= weights[2769];
				12'd2770	: data1 <= weights[2770];
				12'd2771	: data1 <= weights[2771];
				12'd2772	: data1 <= weights[2772];
				12'd2773	: data1 <= weights[2773];
				12'd2774	: data1 <= weights[2774];
				12'd2775	: data1 <= weights[2775];
				12'd2776	: data1 <= weights[2776];
				12'd2777	: data1 <= weights[2777];
				12'd2778	: data1 <= weights[2778];
				12'd2779	: data1 <= weights[2779];
				12'd2780	: data1 <= weights[2780];
				12'd2781	: data1 <= weights[2781];
				12'd2782	: data1 <= weights[2782];
				12'd2783	: data1 <= weights[2783];
				12'd2784	: data1 <= weights[2784];
				12'd2785	: data1 <= weights[2785];
				12'd2786	: data1 <= weights[2786];
				12'd2787	: data1 <= weights[2787];
				12'd2788	: data1 <= weights[2788];
				12'd2789	: data1 <= weights[2789];
				12'd2790	: data1 <= weights[2790];
				12'd2791	: data1 <= weights[2791];
				12'd2792	: data1 <= weights[2792];
				12'd2793	: data1 <= weights[2793];
				12'd2794	: data1 <= weights[2794];
				12'd2795	: data1 <= weights[2795];
				12'd2796	: data1 <= weights[2796];
				12'd2797	: data1 <= weights[2797];
				12'd2798	: data1 <= weights[2798];
				12'd2799	: data1 <= weights[2799];
				12'd2800	: data1 <= weights[2800];
				12'd2801	: data1 <= weights[2801];
				12'd2802	: data1 <= weights[2802];
				12'd2803	: data1 <= weights[2803];
				12'd2804	: data1 <= weights[2804];
				12'd2805	: data1 <= weights[2805];
				12'd2806	: data1 <= weights[2806];
				12'd2807	: data1 <= weights[2807];
				12'd2808	: data1 <= weights[2808];
				12'd2809	: data1 <= weights[2809];
				12'd2810	: data1 <= weights[2810];
				12'd2811	: data1 <= weights[2811];
				12'd2812	: data1 <= weights[2812];
				12'd2813	: data1 <= weights[2813];
				12'd2814	: data1 <= weights[2814];
				12'd2815	: data1 <= weights[2815];
				12'd2816	: data1 <= weights[2816];
				12'd2817	: data1 <= weights[2817];
				12'd2818	: data1 <= weights[2818];
				12'd2819	: data1 <= weights[2819];
				12'd2820	: data1 <= weights[2820];
				12'd2821	: data1 <= weights[2821];
				12'd2822	: data1 <= weights[2822];
				12'd2823	: data1 <= weights[2823];
				12'd2824	: data1 <= weights[2824];
				12'd2825	: data1 <= weights[2825];
				12'd2826	: data1 <= weights[2826];
				12'd2827	: data1 <= weights[2827];
				12'd2828	: data1 <= weights[2828];
				12'd2829	: data1 <= weights[2829];
				12'd2830	: data1 <= weights[2830];
				12'd2831	: data1 <= weights[2831];
				12'd2832	: data1 <= weights[2832];
				12'd2833	: data1 <= weights[2833];
				12'd2834	: data1 <= weights[2834];
				12'd2835	: data1 <= weights[2835];
				12'd2836	: data1 <= weights[2836];
				12'd2837	: data1 <= weights[2837];
				12'd2838	: data1 <= weights[2838];
				12'd2839	: data1 <= weights[2839];
				12'd2840	: data1 <= weights[2840];
				12'd2841	: data1 <= weights[2841];
				12'd2842	: data1 <= weights[2842];
				12'd2843	: data1 <= weights[2843];
				12'd2844	: data1 <= weights[2844];
				12'd2845	: data1 <= weights[2845];
				12'd2846	: data1 <= weights[2846];
				12'd2847	: data1 <= weights[2847];
				12'd2848	: data1 <= weights[2848];
				12'd2849	: data1 <= weights[2849];
				12'd2850	: data1 <= weights[2850];
				12'd2851	: data1 <= weights[2851];
				12'd2852	: data1 <= weights[2852];
				12'd2853	: data1 <= weights[2853];
				12'd2854	: data1 <= weights[2854];
				12'd2855	: data1 <= weights[2855];
				12'd2856	: data1 <= weights[2856];
				12'd2857	: data1 <= weights[2857];
				12'd2858	: data1 <= weights[2858];
				12'd2859	: data1 <= weights[2859];
				12'd2860	: data1 <= weights[2860];
				12'd2861	: data1 <= weights[2861];
				12'd2862	: data1 <= weights[2862];
				12'd2863	: data1 <= weights[2863];
				12'd2864	: data1 <= weights[2864];
				12'd2865	: data1 <= weights[2865];
				12'd2866	: data1 <= weights[2866];
				12'd2867	: data1 <= weights[2867];
				12'd2868	: data1 <= weights[2868];
				12'd2869	: data1 <= weights[2869];
				12'd2870	: data1 <= weights[2870];
				12'd2871	: data1 <= weights[2871];
				12'd2872	: data1 <= weights[2872];
				12'd2873	: data1 <= weights[2873];
				12'd2874	: data1 <= weights[2874];
				12'd2875	: data1 <= weights[2875];
				12'd2876	: data1 <= weights[2876];
				12'd2877	: data1 <= weights[2877];
				12'd2878	: data1 <= weights[2878];
				12'd2879	: data1 <= weights[2879];
				12'd2880	: data1 <= weights[2880];
				12'd2881	: data1 <= weights[2881];
				12'd2882	: data1 <= weights[2882];
				12'd2883	: data1 <= weights[2883];
				12'd2884	: data1 <= weights[2884];
				12'd2885	: data1 <= weights[2885];
				12'd2886	: data1 <= weights[2886];
				12'd2887	: data1 <= weights[2887];
				12'd2888	: data1 <= weights[2888];
				12'd2889	: data1 <= weights[2889];
				12'd2890	: data1 <= weights[2890];
				12'd2891	: data1 <= weights[2891];
				12'd2892	: data1 <= weights[2892];
				12'd2893	: data1 <= weights[2893];
				12'd2894	: data1 <= weights[2894];
				12'd2895	: data1 <= weights[2895];
				12'd2896	: data1 <= weights[2896];
				12'd2897	: data1 <= weights[2897];
				12'd2898	: data1 <= weights[2898];
				12'd2899	: data1 <= weights[2899];
				12'd2900	: data1 <= weights[2900];
				12'd2901	: data1 <= weights[2901];
				12'd2902	: data1 <= weights[2902];
				12'd2903	: data1 <= weights[2903];
				12'd2904	: data1 <= weights[2904];
				12'd2905	: data1 <= weights[2905];
				12'd2906	: data1 <= weights[2906];
				12'd2907	: data1 <= weights[2907];
				12'd2908	: data1 <= weights[2908];
				12'd2909	: data1 <= weights[2909];
				12'd2910	: data1 <= weights[2910];
				12'd2911	: data1 <= weights[2911];
				12'd2912	: data1 <= weights[2912];
				12'd2913	: data1 <= weights[2913];
				12'd2914	: data1 <= weights[2914];
				12'd2915	: data1 <= weights[2915];
				12'd2916	: data1 <= weights[2916];
				12'd2917	: data1 <= weights[2917];
				12'd2918	: data1 <= weights[2918];
				12'd2919	: data1 <= weights[2919];
				12'd2920	: data1 <= weights[2920];
				12'd2921	: data1 <= weights[2921];
				12'd2922	: data1 <= weights[2922];
				12'd2923	: data1 <= weights[2923];
				12'd2924	: data1 <= weights[2924];
				12'd2925	: data1 <= weights[2925];
				12'd2926	: data1 <= weights[2926];
				12'd2927	: data1 <= weights[2927];
				12'd2928	: data1 <= weights[2928];
				12'd2929	: data1 <= weights[2929];
				12'd2930	: data1 <= weights[2930];
				12'd2931	: data1 <= weights[2931];
				12'd2932	: data1 <= weights[2932];
				12'd2933	: data1 <= weights[2933];
				12'd2934	: data1 <= weights[2934];
				12'd2935	: data1 <= weights[2935];
				12'd2936	: data1 <= weights[2936];
				12'd2937	: data1 <= weights[2937];
				12'd2938	: data1 <= weights[2938];
				12'd2939	: data1 <= weights[2939];
				12'd2940	: data1 <= weights[2940];
				12'd2941	: data1 <= weights[2941];
				12'd2942	: data1 <= weights[2942];
				12'd2943	: data1 <= weights[2943];
				12'd2944	: data1 <= weights[2944];
				12'd2945	: data1 <= weights[2945];
				12'd2946	: data1 <= weights[2946];
				12'd2947	: data1 <= weights[2947];
				12'd2948	: data1 <= weights[2948];
				12'd2949	: data1 <= weights[2949];
				12'd2950	: data1 <= weights[2950];
				12'd2951	: data1 <= weights[2951];
				12'd2952	: data1 <= weights[2952];
				12'd2953	: data1 <= weights[2953];
				12'd2954	: data1 <= weights[2954];
				12'd2955	: data1 <= weights[2955];
				12'd2956	: data1 <= weights[2956];
				12'd2957	: data1 <= weights[2957];
				12'd2958	: data1 <= weights[2958];
				12'd2959	: data1 <= weights[2959];
				12'd2960	: data1 <= weights[2960];
				12'd2961	: data1 <= weights[2961];
				12'd2962	: data1 <= weights[2962];
				12'd2963	: data1 <= weights[2963];
				12'd2964	: data1 <= weights[2964];
				12'd2965	: data1 <= weights[2965];
				12'd2966	: data1 <= weights[2966];
				12'd2967	: data1 <= weights[2967];
				12'd2968	: data1 <= weights[2968];
				12'd2969	: data1 <= weights[2969];
				12'd2970	: data1 <= weights[2970];
				12'd2971	: data1 <= weights[2971];
				12'd2972	: data1 <= weights[2972];
				12'd2973	: data1 <= weights[2973];
				12'd2974	: data1 <= weights[2974];
				12'd2975	: data1 <= weights[2975];
				12'd2976	: data1 <= weights[2976];
				12'd2977	: data1 <= weights[2977];
				12'd2978	: data1 <= weights[2978];
				12'd2979	: data1 <= weights[2979];
				12'd2980	: data1 <= weights[2980];
				12'd2981	: data1 <= weights[2981];
				12'd2982	: data1 <= weights[2982];
				12'd2983	: data1 <= weights[2983];
				12'd2984	: data1 <= weights[2984];
				12'd2985	: data1 <= weights[2985];
				12'd2986	: data1 <= weights[2986];
				12'd2987	: data1 <= weights[2987];
				12'd2988	: data1 <= weights[2988];
				12'd2989	: data1 <= weights[2989];
				12'd2990	: data1 <= weights[2990];
				12'd2991	: data1 <= weights[2991];
				12'd2992	: data1 <= weights[2992];
				12'd2993	: data1 <= weights[2993];
				12'd2994	: data1 <= weights[2994];
				12'd2995	: data1 <= weights[2995];
				12'd2996	: data1 <= weights[2996];
				12'd2997	: data1 <= weights[2997];
				12'd2998	: data1 <= weights[2998];
				12'd2999	: data1 <= weights[2999];
				12'd3000	: data1 <= weights[3000];
				12'd3001	: data1 <= weights[3001];
				12'd3002	: data1 <= weights[3002];
				12'd3003	: data1 <= weights[3003];
				12'd3004	: data1 <= weights[3004];
				12'd3005	: data1 <= weights[3005];
				12'd3006	: data1 <= weights[3006];
				12'd3007	: data1 <= weights[3007];
				12'd3008	: data1 <= weights[3008];
				12'd3009	: data1 <= weights[3009];
				12'd3010	: data1 <= weights[3010];
				12'd3011	: data1 <= weights[3011];
				12'd3012	: data1 <= weights[3012];
				12'd3013	: data1 <= weights[3013];
				12'd3014	: data1 <= weights[3014];
				12'd3015	: data1 <= weights[3015];
				12'd3016	: data1 <= weights[3016];
				12'd3017	: data1 <= weights[3017];
				12'd3018	: data1 <= weights[3018];
				12'd3019	: data1 <= weights[3019];
				12'd3020	: data1 <= weights[3020];
				12'd3021	: data1 <= weights[3021];
				12'd3022	: data1 <= weights[3022];
				12'd3023	: data1 <= weights[3023];
				12'd3024	: data1 <= weights[3024];
				12'd3025	: data1 <= weights[3025];
				12'd3026	: data1 <= weights[3026];
				12'd3027	: data1 <= weights[3027];
				12'd3028	: data1 <= weights[3028];
				12'd3029	: data1 <= weights[3029];
				12'd3030	: data1 <= weights[3030];
				12'd3031	: data1 <= weights[3031];
				12'd3032	: data1 <= weights[3032];
				12'd3033	: data1 <= weights[3033];
				12'd3034	: data1 <= weights[3034];
				12'd3035	: data1 <= weights[3035];
				12'd3036	: data1 <= weights[3036];
				12'd3037	: data1 <= weights[3037];
				12'd3038	: data1 <= weights[3038];
				12'd3039	: data1 <= weights[3039];
				12'd3040	: data1 <= weights[3040];
				12'd3041	: data1 <= weights[3041];
				12'd3042	: data1 <= weights[3042];
				12'd3043	: data1 <= weights[3043];
				12'd3044	: data1 <= weights[3044];
				12'd3045	: data1 <= weights[3045];
				12'd3046	: data1 <= weights[3046];
				12'd3047	: data1 <= weights[3047];
				12'd3048	: data1 <= weights[3048];
				12'd3049	: data1 <= weights[3049];
				12'd3050	: data1 <= weights[3050];
				12'd3051	: data1 <= weights[3051];
				12'd3052	: data1 <= weights[3052];
				12'd3053	: data1 <= weights[3053];
				12'd3054	: data1 <= weights[3054];
				12'd3055	: data1 <= weights[3055];
				12'd3056	: data1 <= weights[3056];
				12'd3057	: data1 <= weights[3057];
				12'd3058	: data1 <= weights[3058];
				12'd3059	: data1 <= weights[3059];
				12'd3060	: data1 <= weights[3060];
				12'd3061	: data1 <= weights[3061];
				12'd3062	: data1 <= weights[3062];
				12'd3063	: data1 <= weights[3063];
				12'd3064	: data1 <= weights[3064];
				12'd3065	: data1 <= weights[3065];
				12'd3066	: data1 <= weights[3066];
				12'd3067	: data1 <= weights[3067];
				12'd3068	: data1 <= weights[3068];
				12'd3069	: data1 <= weights[3069];
				12'd3070	: data1 <= weights[3070];
				12'd3071	: data1 <= weights[3071];
				12'd3072	: data1 <= weights[3072];
				12'd3073	: data1 <= weights[3073];
				12'd3074	: data1 <= weights[3074];
				12'd3075	: data1 <= weights[3075];
				12'd3076	: data1 <= weights[3076];
				12'd3077	: data1 <= weights[3077];
				12'd3078	: data1 <= weights[3078];
				12'd3079	: data1 <= weights[3079];
				12'd3080	: data1 <= weights[3080];
				12'd3081	: data1 <= weights[3081];
				12'd3082	: data1 <= weights[3082];
				12'd3083	: data1 <= weights[3083];
				12'd3084	: data1 <= weights[3084];
				12'd3085	: data1 <= weights[3085];
				12'd3086	: data1 <= weights[3086];
				12'd3087	: data1 <= weights[3087];
				12'd3088	: data1 <= weights[3088];
				12'd3089	: data1 <= weights[3089];
				12'd3090	: data1 <= weights[3090];
				12'd3091	: data1 <= weights[3091];
				12'd3092	: data1 <= weights[3092];
				12'd3093	: data1 <= weights[3093];
				12'd3094	: data1 <= weights[3094];
				12'd3095	: data1 <= weights[3095];
				12'd3096	: data1 <= weights[3096];
				12'd3097	: data1 <= weights[3097];
				12'd3098	: data1 <= weights[3098];
				12'd3099	: data1 <= weights[3099];
				12'd3100	: data1 <= weights[3100];
				12'd3101	: data1 <= weights[3101];
				12'd3102	: data1 <= weights[3102];
				12'd3103	: data1 <= weights[3103];
				12'd3104	: data1 <= weights[3104];
				12'd3105	: data1 <= weights[3105];
				12'd3106	: data1 <= weights[3106];
				12'd3107	: data1 <= weights[3107];
				12'd3108	: data1 <= weights[3108];
				12'd3109	: data1 <= weights[3109];
				12'd3110	: data1 <= weights[3110];
				12'd3111	: data1 <= weights[3111];
				12'd3112	: data1 <= weights[3112];
				12'd3113	: data1 <= weights[3113];
				12'd3114	: data1 <= weights[3114];
				12'd3115	: data1 <= weights[3115];
				12'd3116	: data1 <= weights[3116];
				12'd3117	: data1 <= weights[3117];
				12'd3118	: data1 <= weights[3118];
				12'd3119	: data1 <= weights[3119];
				12'd3120	: data1 <= weights[3120];
				12'd3121	: data1 <= weights[3121];
				12'd3122	: data1 <= weights[3122];
				12'd3123	: data1 <= weights[3123];
				12'd3124	: data1 <= weights[3124];
				12'd3125	: data1 <= weights[3125];
				12'd3126	: data1 <= weights[3126];
				12'd3127	: data1 <= weights[3127];
				12'd3128	: data1 <= weights[3128];
				12'd3129	: data1 <= weights[3129];
				12'd3130	: data1 <= weights[3130];
				12'd3131	: data1 <= weights[3131];
				12'd3132	: data1 <= weights[3132];
				12'd3133	: data1 <= weights[3133];
				12'd3134	: data1 <= weights[3134];
				12'd3135	: data1 <= weights[3135];
				12'd3136	: data1 <= weights[3136];
				12'd3137	: data1 <= weights[3137];
				12'd3138	: data1 <= weights[3138];
				12'd3139	: data1 <= weights[3139];
				12'd3140	: data1 <= weights[3140];
				12'd3141	: data1 <= weights[3141];
				12'd3142	: data1 <= weights[3142];
				12'd3143	: data1 <= weights[3143];
				12'd3144	: data1 <= weights[3144];
				12'd3145	: data1 <= weights[3145];
				12'd3146	: data1 <= weights[3146];
				12'd3147	: data1 <= weights[3147];
				12'd3148	: data1 <= weights[3148];
				12'd3149	: data1 <= weights[3149];
				12'd3150	: data1 <= weights[3150];
				12'd3151	: data1 <= weights[3151];
				12'd3152	: data1 <= weights[3152];
				12'd3153	: data1 <= weights[3153];
				12'd3154	: data1 <= weights[3154];
				12'd3155	: data1 <= weights[3155];
				12'd3156	: data1 <= weights[3156];
				12'd3157	: data1 <= weights[3157];
				12'd3158	: data1 <= weights[3158];
				12'd3159	: data1 <= weights[3159];
				12'd3160	: data1 <= weights[3160];
				12'd3161	: data1 <= weights[3161];
				12'd3162	: data1 <= weights[3162];
				12'd3163	: data1 <= weights[3163];
				12'd3164	: data1 <= weights[3164];
				12'd3165	: data1 <= weights[3165];
				12'd3166	: data1 <= weights[3166];
				12'd3167	: data1 <= weights[3167];
				12'd3168	: data1 <= weights[3168];
				12'd3169	: data1 <= weights[3169];
				12'd3170	: data1 <= weights[3170];
				12'd3171	: data1 <= weights[3171];
				12'd3172	: data1 <= weights[3172];
				12'd3173	: data1 <= weights[3173];
				12'd3174	: data1 <= weights[3174];
				12'd3175	: data1 <= weights[3175];
				12'd3176	: data1 <= weights[3176];
				12'd3177	: data1 <= weights[3177];
				12'd3178	: data1 <= weights[3178];
				12'd3179	: data1 <= weights[3179];
				12'd3180	: data1 <= weights[3180];
				12'd3181	: data1 <= weights[3181];
				12'd3182	: data1 <= weights[3182];
				12'd3183	: data1 <= weights[3183];
				12'd3184	: data1 <= weights[3184];
				12'd3185	: data1 <= weights[3185];
				12'd3186	: data1 <= weights[3186];
				12'd3187	: data1 <= weights[3187];
				12'd3188	: data1 <= weights[3188];
				12'd3189	: data1 <= weights[3189];
				12'd3190	: data1 <= weights[3190];
				12'd3191	: data1 <= weights[3191];
				12'd3192	: data1 <= weights[3192];
				12'd3193	: data1 <= weights[3193];
				12'd3194	: data1 <= weights[3194];
				12'd3195	: data1 <= weights[3195];
				12'd3196	: data1 <= weights[3196];
				12'd3197	: data1 <= weights[3197];
				12'd3198	: data1 <= weights[3198];
				12'd3199	: data1 <= weights[3199];
				12'd3200	: data1 <= weights[3200];
				12'd3201	: data1 <= weights[3201];
				12'd3202	: data1 <= weights[3202];
				12'd3203	: data1 <= weights[3203];
				12'd3204	: data1 <= weights[3204];
				12'd3205	: data1 <= weights[3205];
				12'd3206	: data1 <= weights[3206];
				12'd3207	: data1 <= weights[3207];
				12'd3208	: data1 <= weights[3208];
				12'd3209	: data1 <= weights[3209];
				12'd3210	: data1 <= weights[3210];
				12'd3211	: data1 <= weights[3211];
				12'd3212	: data1 <= weights[3212];
				12'd3213	: data1 <= weights[3213];
				12'd3214	: data1 <= weights[3214];
				12'd3215	: data1 <= weights[3215];
				12'd3216	: data1 <= weights[3216];
				12'd3217	: data1 <= weights[3217];
				12'd3218	: data1 <= weights[3218];
				12'd3219	: data1 <= weights[3219];
				12'd3220	: data1 <= weights[3220];
				12'd3221	: data1 <= weights[3221];
				12'd3222	: data1 <= weights[3222];
				12'd3223	: data1 <= weights[3223];
				12'd3224	: data1 <= weights[3224];
				12'd3225	: data1 <= weights[3225];
				12'd3226	: data1 <= weights[3226];
				12'd3227	: data1 <= weights[3227];
				12'd3228	: data1 <= weights[3228];
				12'd3229	: data1 <= weights[3229];
				12'd3230	: data1 <= weights[3230];
				12'd3231	: data1 <= weights[3231];
				12'd3232	: data1 <= weights[3232];
				12'd3233	: data1 <= weights[3233];
				12'd3234	: data1 <= weights[3234];
				12'd3235	: data1 <= weights[3235];
				12'd3236	: data1 <= weights[3236];
				12'd3237	: data1 <= weights[3237];
				12'd3238	: data1 <= weights[3238];
				12'd3239	: data1 <= weights[3239];
				12'd3240	: data1 <= weights[3240];
				12'd3241	: data1 <= weights[3241];
				12'd3242	: data1 <= weights[3242];
				12'd3243	: data1 <= weights[3243];
				12'd3244	: data1 <= weights[3244];
				12'd3245	: data1 <= weights[3245];
				12'd3246	: data1 <= weights[3246];
				12'd3247	: data1 <= weights[3247];
				12'd3248	: data1 <= weights[3248];
				12'd3249	: data1 <= weights[3249];
				12'd3250	: data1 <= weights[3250];
				12'd3251	: data1 <= weights[3251];
				12'd3252	: data1 <= weights[3252];
				12'd3253	: data1 <= weights[3253];
				12'd3254	: data1 <= weights[3254];
				12'd3255	: data1 <= weights[3255];
				12'd3256	: data1 <= weights[3256];
				12'd3257	: data1 <= weights[3257];
				12'd3258	: data1 <= weights[3258];
				12'd3259	: data1 <= weights[3259];
				12'd3260	: data1 <= weights[3260];
				12'd3261	: data1 <= weights[3261];
				12'd3262	: data1 <= weights[3262];
				12'd3263	: data1 <= weights[3263];
				12'd3264	: data1 <= weights[3264];
				12'd3265	: data1 <= weights[3265];
				12'd3266	: data1 <= weights[3266];
				12'd3267	: data1 <= weights[3267];
				12'd3268	: data1 <= weights[3268];
				12'd3269	: data1 <= weights[3269];
				12'd3270	: data1 <= weights[3270];
				12'd3271	: data1 <= weights[3271];
				12'd3272	: data1 <= weights[3272];
				12'd3273	: data1 <= weights[3273];
				12'd3274	: data1 <= weights[3274];
				12'd3275	: data1 <= weights[3275];
				12'd3276	: data1 <= weights[3276];
				12'd3277	: data1 <= weights[3277];
				12'd3278	: data1 <= weights[3278];
				12'd3279	: data1 <= weights[3279];
				12'd3280	: data1 <= weights[3280];
				12'd3281	: data1 <= weights[3281];
				12'd3282	: data1 <= weights[3282];
				12'd3283	: data1 <= weights[3283];
				12'd3284	: data1 <= weights[3284];
				12'd3285	: data1 <= weights[3285];
				12'd3286	: data1 <= weights[3286];
				12'd3287	: data1 <= weights[3287];
				12'd3288	: data1 <= weights[3288];
				12'd3289	: data1 <= weights[3289];
				12'd3290	: data1 <= weights[3290];
				12'd3291	: data1 <= weights[3291];
				12'd3292	: data1 <= weights[3292];
				12'd3293	: data1 <= weights[3293];
				12'd3294	: data1 <= weights[3294];
				12'd3295	: data1 <= weights[3295];
				12'd3296	: data1 <= weights[3296];
				12'd3297	: data1 <= weights[3297];
				12'd3298	: data1 <= weights[3298];
				12'd3299	: data1 <= weights[3299];
				12'd3300	: data1 <= weights[3300];
				12'd3301	: data1 <= weights[3301];
				12'd3302	: data1 <= weights[3302];
				12'd3303	: data1 <= weights[3303];
				12'd3304	: data1 <= weights[3304];
				12'd3305	: data1 <= weights[3305];
				12'd3306	: data1 <= weights[3306];
				12'd3307	: data1 <= weights[3307];
				12'd3308	: data1 <= weights[3308];
				12'd3309	: data1 <= weights[3309];
				12'd3310	: data1 <= weights[3310];
				12'd3311	: data1 <= weights[3311];
				12'd3312	: data1 <= weights[3312];
				12'd3313	: data1 <= weights[3313];
				12'd3314	: data1 <= weights[3314];
				12'd3315	: data1 <= weights[3315];
				12'd3316	: data1 <= weights[3316];
				12'd3317	: data1 <= weights[3317];
				12'd3318	: data1 <= weights[3318];
				12'd3319	: data1 <= weights[3319];
				12'd3320	: data1 <= weights[3320];
				12'd3321	: data1 <= weights[3321];
				12'd3322	: data1 <= weights[3322];
				12'd3323	: data1 <= weights[3323];
				12'd3324	: data1 <= weights[3324];
				12'd3325	: data1 <= weights[3325];
				12'd3326	: data1 <= weights[3326];
				12'd3327	: data1 <= weights[3327];
				12'd3328	: data1 <= weights[3328];
				12'd3329	: data1 <= weights[3329];
				12'd3330	: data1 <= weights[3330];
				12'd3331	: data1 <= weights[3331];
				12'd3332	: data1 <= weights[3332];
				12'd3333	: data1 <= weights[3333];
				12'd3334	: data1 <= weights[3334];
				12'd3335	: data1 <= weights[3335];
				12'd3336	: data1 <= weights[3336];
				12'd3337	: data1 <= weights[3337];
				12'd3338	: data1 <= weights[3338];
				12'd3339	: data1 <= weights[3339];
				12'd3340	: data1 <= weights[3340];
				12'd3341	: data1 <= weights[3341];
				12'd3342	: data1 <= weights[3342];
				12'd3343	: data1 <= weights[3343];
				12'd3344	: data1 <= weights[3344];
				12'd3345	: data1 <= weights[3345];
				12'd3346	: data1 <= weights[3346];
				12'd3347	: data1 <= weights[3347];
				12'd3348	: data1 <= weights[3348];
				12'd3349	: data1 <= weights[3349];
				12'd3350	: data1 <= weights[3350];
				12'd3351	: data1 <= weights[3351];
				12'd3352	: data1 <= weights[3352];
				12'd3353	: data1 <= weights[3353];
				12'd3354	: data1 <= weights[3354];
				12'd3355	: data1 <= weights[3355];
				12'd3356	: data1 <= weights[3356];
				12'd3357	: data1 <= weights[3357];
				12'd3358	: data1 <= weights[3358];
				12'd3359	: data1 <= weights[3359];
				12'd3360	: data1 <= weights[3360];
				12'd3361	: data1 <= weights[3361];
				12'd3362	: data1 <= weights[3362];
				12'd3363	: data1 <= weights[3363];
				12'd3364	: data1 <= weights[3364];
				12'd3365	: data1 <= weights[3365];
				12'd3366	: data1 <= weights[3366];
				12'd3367	: data1 <= weights[3367];
				12'd3368	: data1 <= weights[3368];
				12'd3369	: data1 <= weights[3369];
				12'd3370	: data1 <= weights[3370];
				12'd3371	: data1 <= weights[3371];
				12'd3372	: data1 <= weights[3372];
				12'd3373	: data1 <= weights[3373];
				12'd3374	: data1 <= weights[3374];
				12'd3375	: data1 <= weights[3375];
				12'd3376	: data1 <= weights[3376];
				12'd3377	: data1 <= weights[3377];
				12'd3378	: data1 <= weights[3378];
				12'd3379	: data1 <= weights[3379];
				12'd3380	: data1 <= weights[3380];
				12'd3381	: data1 <= weights[3381];
				12'd3382	: data1 <= weights[3382];
				12'd3383	: data1 <= weights[3383];
				12'd3384	: data1 <= weights[3384];
				12'd3385	: data1 <= weights[3385];
				12'd3386	: data1 <= weights[3386];
				12'd3387	: data1 <= weights[3387];
				12'd3388	: data1 <= weights[3388];
				12'd3389	: data1 <= weights[3389];
				12'd3390	: data1 <= weights[3390];
				12'd3391	: data1 <= weights[3391];
				12'd3392	: data1 <= weights[3392];
				12'd3393	: data1 <= weights[3393];
				12'd3394	: data1 <= weights[3394];
				12'd3395	: data1 <= weights[3395];
				12'd3396	: data1 <= weights[3396];
				12'd3397	: data1 <= weights[3397];
				12'd3398	: data1 <= weights[3398];
				12'd3399	: data1 <= weights[3399];
				12'd3400	: data1 <= weights[3400];
				12'd3401	: data1 <= weights[3401];
				12'd3402	: data1 <= weights[3402];
				12'd3403	: data1 <= weights[3403];
				12'd3404	: data1 <= weights[3404];
				12'd3405	: data1 <= weights[3405];
				12'd3406	: data1 <= weights[3406];
				12'd3407	: data1 <= weights[3407];
				12'd3408	: data1 <= weights[3408];
				12'd3409	: data1 <= weights[3409];
				12'd3410	: data1 <= weights[3410];
				12'd3411	: data1 <= weights[3411];
				12'd3412	: data1 <= weights[3412];
				12'd3413	: data1 <= weights[3413];
				12'd3414	: data1 <= weights[3414];
				12'd3415	: data1 <= weights[3415];
				12'd3416	: data1 <= weights[3416];
				12'd3417	: data1 <= weights[3417];
				12'd3418	: data1 <= weights[3418];
				12'd3419	: data1 <= weights[3419];
				12'd3420	: data1 <= weights[3420];
				12'd3421	: data1 <= weights[3421];
				12'd3422	: data1 <= weights[3422];
				12'd3423	: data1 <= weights[3423];
				12'd3424	: data1 <= weights[3424];
				12'd3425	: data1 <= weights[3425];
				12'd3426	: data1 <= weights[3426];
				12'd3427	: data1 <= weights[3427];
				12'd3428	: data1 <= weights[3428];
				12'd3429	: data1 <= weights[3429];
				12'd3430	: data1 <= weights[3430];
				12'd3431	: data1 <= weights[3431];
				12'd3432	: data1 <= weights[3432];
				12'd3433	: data1 <= weights[3433];
				12'd3434	: data1 <= weights[3434];
				12'd3435	: data1 <= weights[3435];
				12'd3436	: data1 <= weights[3436];
				12'd3437	: data1 <= weights[3437];
				12'd3438	: data1 <= weights[3438];
				12'd3439	: data1 <= weights[3439];
				12'd3440	: data1 <= weights[3440];
				12'd3441	: data1 <= weights[3441];
				12'd3442	: data1 <= weights[3442];
				12'd3443	: data1 <= weights[3443];
				12'd3444	: data1 <= weights[3444];
				12'd3445	: data1 <= weights[3445];
				12'd3446	: data1 <= weights[3446];
				12'd3447	: data1 <= weights[3447];
				12'd3448	: data1 <= weights[3448];
				12'd3449	: data1 <= weights[3449];
				12'd3450	: data1 <= weights[3450];
				12'd3451	: data1 <= weights[3451];
				12'd3452	: data1 <= weights[3452];
				12'd3453	: data1 <= weights[3453];
				12'd3454	: data1 <= weights[3454];
				12'd3455	: data1 <= weights[3455];
				12'd3456	: data1 <= weights[3456];
				12'd3457	: data1 <= weights[3457];
				12'd3458	: data1 <= weights[3458];
				12'd3459	: data1 <= weights[3459];
				12'd3460	: data1 <= weights[3460];
				12'd3461	: data1 <= weights[3461];
				12'd3462	: data1 <= weights[3462];
				12'd3463	: data1 <= weights[3463];
				12'd3464	: data1 <= weights[3464];
				12'd3465	: data1 <= weights[3465];
				12'd3466	: data1 <= weights[3466];
				12'd3467	: data1 <= weights[3467];
				12'd3468	: data1 <= weights[3468];
				12'd3469	: data1 <= weights[3469];
				12'd3470	: data1 <= weights[3470];
				12'd3471	: data1 <= weights[3471];
				12'd3472	: data1 <= weights[3472];
				12'd3473	: data1 <= weights[3473];
				12'd3474	: data1 <= weights[3474];
				12'd3475	: data1 <= weights[3475];
				12'd3476	: data1 <= weights[3476];
				12'd3477	: data1 <= weights[3477];
				12'd3478	: data1 <= weights[3478];
				12'd3479	: data1 <= weights[3479];
				12'd3480	: data1 <= weights[3480];
				12'd3481	: data1 <= weights[3481];
				12'd3482	: data1 <= weights[3482];
				12'd3483	: data1 <= weights[3483];
				12'd3484	: data1 <= weights[3484];
				12'd3485	: data1 <= weights[3485];
				12'd3486	: data1 <= weights[3486];
				12'd3487	: data1 <= weights[3487];
				12'd3488	: data1 <= weights[3488];
				12'd3489	: data1 <= weights[3489];
				12'd3490	: data1 <= weights[3490];
				12'd3491	: data1 <= weights[3491];
				12'd3492	: data1 <= weights[3492];
				12'd3493	: data1 <= weights[3493];
				12'd3494	: data1 <= weights[3494];
				12'd3495	: data1 <= weights[3495];
				12'd3496	: data1 <= weights[3496];
				12'd3497	: data1 <= weights[3497];
				12'd3498	: data1 <= weights[3498];
				12'd3499	: data1 <= weights[3499];
				12'd3500	: data1 <= weights[3500];
				12'd3501	: data1 <= weights[3501];
				12'd3502	: data1 <= weights[3502];
				12'd3503	: data1 <= weights[3503];
				12'd3504	: data1 <= weights[3504];
				12'd3505	: data1 <= weights[3505];
				12'd3506	: data1 <= weights[3506];
				12'd3507	: data1 <= weights[3507];
				12'd3508	: data1 <= weights[3508];
				12'd3509	: data1 <= weights[3509];
				12'd3510	: data1 <= weights[3510];
				12'd3511	: data1 <= weights[3511];
				12'd3512	: data1 <= weights[3512];
				12'd3513	: data1 <= weights[3513];
				12'd3514	: data1 <= weights[3514];
				12'd3515	: data1 <= weights[3515];
				12'd3516	: data1 <= weights[3516];
				12'd3517	: data1 <= weights[3517];
				12'd3518	: data1 <= weights[3518];
				12'd3519	: data1 <= weights[3519];
				12'd3520	: data1 <= weights[3520];
				12'd3521	: data1 <= weights[3521];
				12'd3522	: data1 <= weights[3522];
				12'd3523	: data1 <= weights[3523];
				12'd3524	: data1 <= weights[3524];
				12'd3525	: data1 <= weights[3525];
				12'd3526	: data1 <= weights[3526];
				12'd3527	: data1 <= weights[3527];
				12'd3528	: data1 <= weights[3528];
				12'd3529	: data1 <= weights[3529];
				12'd3530	: data1 <= weights[3530];
				12'd3531	: data1 <= weights[3531];
				12'd3532	: data1 <= weights[3532];
				12'd3533	: data1 <= weights[3533];
				12'd3534	: data1 <= weights[3534];
				12'd3535	: data1 <= weights[3535];
				12'd3536	: data1 <= weights[3536];
				12'd3537	: data1 <= weights[3537];
				12'd3538	: data1 <= weights[3538];
				12'd3539	: data1 <= weights[3539];
				12'd3540	: data1 <= weights[3540];
				12'd3541	: data1 <= weights[3541];
				12'd3542	: data1 <= weights[3542];
				12'd3543	: data1 <= weights[3543];
				12'd3544	: data1 <= weights[3544];
				12'd3545	: data1 <= weights[3545];
				12'd3546	: data1 <= weights[3546];
				12'd3547	: data1 <= weights[3547];
				12'd3548	: data1 <= weights[3548];
				12'd3549	: data1 <= weights[3549];
				12'd3550	: data1 <= weights[3550];
				12'd3551	: data1 <= weights[3551];
				12'd3552	: data1 <= weights[3552];
				12'd3553	: data1 <= weights[3553];
				12'd3554	: data1 <= weights[3554];
				12'd3555	: data1 <= weights[3555];
				12'd3556	: data1 <= weights[3556];
				12'd3557	: data1 <= weights[3557];
				12'd3558	: data1 <= weights[3558];
				12'd3559	: data1 <= weights[3559];
				12'd3560	: data1 <= weights[3560];
				12'd3561	: data1 <= weights[3561];
				12'd3562	: data1 <= weights[3562];
				12'd3563	: data1 <= weights[3563];
				12'd3564	: data1 <= weights[3564];
				12'd3565	: data1 <= weights[3565];
				12'd3566	: data1 <= weights[3566];
				12'd3567	: data1 <= weights[3567];
				12'd3568	: data1 <= weights[3568];
				12'd3569	: data1 <= weights[3569];
				12'd3570	: data1 <= weights[3570];
				12'd3571	: data1 <= weights[3571];
				12'd3572	: data1 <= weights[3572];
				12'd3573	: data1 <= weights[3573];
				12'd3574	: data1 <= weights[3574];
				12'd3575	: data1 <= weights[3575];
				12'd3576	: data1 <= weights[3576];
				12'd3577	: data1 <= weights[3577];
				12'd3578	: data1 <= weights[3578];
				12'd3579	: data1 <= weights[3579];
				12'd3580	: data1 <= weights[3580];
				12'd3581	: data1 <= weights[3581];
				12'd3582	: data1 <= weights[3582];
				12'd3583	: data1 <= weights[3583];
				12'd3584	: data1 <= weights[3584];
				12'd3585	: data1 <= weights[3585];
				12'd3586	: data1 <= weights[3586];
				12'd3587	: data1 <= weights[3587];
				12'd3588	: data1 <= weights[3588];
				12'd3589	: data1 <= weights[3589];
				12'd3590	: data1 <= weights[3590];
				12'd3591	: data1 <= weights[3591];
				12'd3592	: data1 <= weights[3592];
				12'd3593	: data1 <= weights[3593];
				12'd3594	: data1 <= weights[3594];
				12'd3595	: data1 <= weights[3595];
				12'd3596	: data1 <= weights[3596];
				12'd3597	: data1 <= weights[3597];
				12'd3598	: data1 <= weights[3598];
				12'd3599	: data1 <= weights[3599];
				12'd3600	: data1 <= weights[3600];
				12'd3601	: data1 <= weights[3601];
				12'd3602	: data1 <= weights[3602];
				12'd3603	: data1 <= weights[3603];
				12'd3604	: data1 <= weights[3604];
				12'd3605	: data1 <= weights[3605];
				12'd3606	: data1 <= weights[3606];
				12'd3607	: data1 <= weights[3607];
				12'd3608	: data1 <= weights[3608];
				12'd3609	: data1 <= weights[3609];
				12'd3610	: data1 <= weights[3610];
				12'd3611	: data1 <= weights[3611];
				12'd3612	: data1 <= weights[3612];
				12'd3613	: data1 <= weights[3613];
				12'd3614	: data1 <= weights[3614];
				12'd3615	: data1 <= weights[3615];
				12'd3616	: data1 <= weights[3616];
				12'd3617	: data1 <= weights[3617];
				12'd3618	: data1 <= weights[3618];
				12'd3619	: data1 <= weights[3619];
				12'd3620	: data1 <= weights[3620];
				12'd3621	: data1 <= weights[3621];
				12'd3622	: data1 <= weights[3622];
				12'd3623	: data1 <= weights[3623];
				12'd3624	: data1 <= weights[3624];
				12'd3625	: data1 <= weights[3625];
				12'd3626	: data1 <= weights[3626];
				12'd3627	: data1 <= weights[3627];
				12'd3628	: data1 <= weights[3628];
				12'd3629	: data1 <= weights[3629];
				12'd3630	: data1 <= weights[3630];
				12'd3631	: data1 <= weights[3631];
				12'd3632	: data1 <= weights[3632];
				12'd3633	: data1 <= weights[3633];
				12'd3634	: data1 <= weights[3634];
				12'd3635	: data1 <= weights[3635];
				12'd3636	: data1 <= weights[3636];
				12'd3637	: data1 <= weights[3637];
				12'd3638	: data1 <= weights[3638];
				12'd3639	: data1 <= weights[3639];
				12'd3640	: data1 <= weights[3640];
				12'd3641	: data1 <= weights[3641];
				12'd3642	: data1 <= weights[3642];
				12'd3643	: data1 <= weights[3643];
				12'd3644	: data1 <= weights[3644];
				12'd3645	: data1 <= weights[3645];
				12'd3646	: data1 <= weights[3646];
				12'd3647	: data1 <= weights[3647];
				12'd3648	: data1 <= weights[3648];
				12'd3649	: data1 <= weights[3649];
				12'd3650	: data1 <= weights[3650];
				12'd3651	: data1 <= weights[3651];
				12'd3652	: data1 <= weights[3652];
				12'd3653	: data1 <= weights[3653];
				12'd3654	: data1 <= weights[3654];
				12'd3655	: data1 <= weights[3655];
				12'd3656	: data1 <= weights[3656];
				12'd3657	: data1 <= weights[3657];
				12'd3658	: data1 <= weights[3658];
				12'd3659	: data1 <= weights[3659];
				12'd3660	: data1 <= weights[3660];
				12'd3661	: data1 <= weights[3661];
				12'd3662	: data1 <= weights[3662];
				12'd3663	: data1 <= weights[3663];
				12'd3664	: data1 <= weights[3664];
				12'd3665	: data1 <= weights[3665];
				12'd3666	: data1 <= weights[3666];
				12'd3667	: data1 <= weights[3667];
				12'd3668	: data1 <= weights[3668];
				12'd3669	: data1 <= weights[3669];
				12'd3670	: data1 <= weights[3670];
				12'd3671	: data1 <= weights[3671];
				12'd3672	: data1 <= weights[3672];
				12'd3673	: data1 <= weights[3673];
				12'd3674	: data1 <= weights[3674];
				12'd3675	: data1 <= weights[3675];
				12'd3676	: data1 <= weights[3676];
				12'd3677	: data1 <= weights[3677];
				12'd3678	: data1 <= weights[3678];
				12'd3679	: data1 <= weights[3679];
				12'd3680	: data1 <= weights[3680];
				12'd3681	: data1 <= weights[3681];
				12'd3682	: data1 <= weights[3682];
				12'd3683	: data1 <= weights[3683];
				12'd3684	: data1 <= weights[3684];
				12'd3685	: data1 <= weights[3685];
				12'd3686	: data1 <= weights[3686];
				12'd3687	: data1 <= weights[3687];
				12'd3688	: data1 <= weights[3688];
				12'd3689	: data1 <= weights[3689];
				12'd3690	: data1 <= weights[3690];
				12'd3691	: data1 <= weights[3691];
				12'd3692	: data1 <= weights[3692];
				12'd3693	: data1 <= weights[3693];
				12'd3694	: data1 <= weights[3694];
				12'd3695	: data1 <= weights[3695];
				12'd3696	: data1 <= weights[3696];
				12'd3697	: data1 <= weights[3697];
				12'd3698	: data1 <= weights[3698];
				12'd3699	: data1 <= weights[3699];
				12'd3700	: data1 <= weights[3700];
				12'd3701	: data1 <= weights[3701];
				12'd3702	: data1 <= weights[3702];
				12'd3703	: data1 <= weights[3703];
				12'd3704	: data1 <= weights[3704];
				12'd3705	: data1 <= weights[3705];
				12'd3706	: data1 <= weights[3706];
				12'd3707	: data1 <= weights[3707];
				12'd3708	: data1 <= weights[3708];
				12'd3709	: data1 <= weights[3709];
				12'd3710	: data1 <= weights[3710];
				12'd3711	: data1 <= weights[3711];
				12'd3712	: data1 <= weights[3712];
				12'd3713	: data1 <= weights[3713];
				12'd3714	: data1 <= weights[3714];
				12'd3715	: data1 <= weights[3715];
				12'd3716	: data1 <= weights[3716];
				12'd3717	: data1 <= weights[3717];
				12'd3718	: data1 <= weights[3718];
				12'd3719	: data1 <= weights[3719];
				12'd3720	: data1 <= weights[3720];
				12'd3721	: data1 <= weights[3721];
				12'd3722	: data1 <= weights[3722];
				12'd3723	: data1 <= weights[3723];
				12'd3724	: data1 <= weights[3724];
				12'd3725	: data1 <= weights[3725];
				12'd3726	: data1 <= weights[3726];
				12'd3727	: data1 <= weights[3727];
				12'd3728	: data1 <= weights[3728];
				12'd3729	: data1 <= weights[3729];
				12'd3730	: data1 <= weights[3730];
				12'd3731	: data1 <= weights[3731];
				12'd3732	: data1 <= weights[3732];
				12'd3733	: data1 <= weights[3733];
				12'd3734	: data1 <= weights[3734];
				12'd3735	: data1 <= weights[3735];
				12'd3736	: data1 <= weights[3736];
				12'd3737	: data1 <= weights[3737];
				12'd3738	: data1 <= weights[3738];
				12'd3739	: data1 <= weights[3739];
				12'd3740	: data1 <= weights[3740];
				12'd3741	: data1 <= weights[3741];
				12'd3742	: data1 <= weights[3742];
				12'd3743	: data1 <= weights[3743];
				12'd3744	: data1 <= weights[3744];
				12'd3745	: data1 <= weights[3745];
				12'd3746	: data1 <= weights[3746];
				12'd3747	: data1 <= weights[3747];
				12'd3748	: data1 <= weights[3748];
				12'd3749	: data1 <= weights[3749];
				12'd3750	: data1 <= weights[3750];
				12'd3751	: data1 <= weights[3751];
				12'd3752	: data1 <= weights[3752];
				12'd3753	: data1 <= weights[3753];
				12'd3754	: data1 <= weights[3754];
				12'd3755	: data1 <= weights[3755];
				12'd3756	: data1 <= weights[3756];
				12'd3757	: data1 <= weights[3757];
				12'd3758	: data1 <= weights[3758];
				12'd3759	: data1 <= weights[3759];
				12'd3760	: data1 <= weights[3760];
				12'd3761	: data1 <= weights[3761];
				12'd3762	: data1 <= weights[3762];
				12'd3763	: data1 <= weights[3763];
				12'd3764	: data1 <= weights[3764];
				12'd3765	: data1 <= weights[3765];
				12'd3766	: data1 <= weights[3766];
				12'd3767	: data1 <= weights[3767];
				12'd3768	: data1 <= weights[3768];
				12'd3769	: data1 <= weights[3769];
				12'd3770	: data1 <= weights[3770];
				12'd3771	: data1 <= weights[3771];
				12'd3772	: data1 <= weights[3772];
				12'd3773	: data1 <= weights[3773];
				12'd3774	: data1 <= weights[3774];
				12'd3775	: data1 <= weights[3775];
				12'd3776	: data1 <= weights[3776];
				12'd3777	: data1 <= weights[3777];
				12'd3778	: data1 <= weights[3778];
				12'd3779	: data1 <= weights[3779];
				12'd3780	: data1 <= weights[3780];
				12'd3781	: data1 <= weights[3781];
				12'd3782	: data1 <= weights[3782];
				12'd3783	: data1 <= weights[3783];
				12'd3784	: data1 <= weights[3784];
				12'd3785	: data1 <= weights[3785];
				12'd3786	: data1 <= weights[3786];
				12'd3787	: data1 <= weights[3787];
				12'd3788	: data1 <= weights[3788];
				12'd3789	: data1 <= weights[3789];
				12'd3790	: data1 <= weights[3790];
				12'd3791	: data1 <= weights[3791];
				12'd3792	: data1 <= weights[3792];
				12'd3793	: data1 <= weights[3793];
				12'd3794	: data1 <= weights[3794];
				12'd3795	: data1 <= weights[3795];
				12'd3796	: data1 <= weights[3796];
				12'd3797	: data1 <= weights[3797];
				12'd3798	: data1 <= weights[3798];
				12'd3799	: data1 <= weights[3799];
				12'd3800	: data1 <= weights[3800];
				12'd3801	: data1 <= weights[3801];
				12'd3802	: data1 <= weights[3802];
				12'd3803	: data1 <= weights[3803];
				12'd3804	: data1 <= weights[3804];
				12'd3805	: data1 <= weights[3805];
				12'd3806	: data1 <= weights[3806];
				12'd3807	: data1 <= weights[3807];
				12'd3808	: data1 <= weights[3808];
				12'd3809	: data1 <= weights[3809];
				12'd3810	: data1 <= weights[3810];
				12'd3811	: data1 <= weights[3811];
				12'd3812	: data1 <= weights[3812];
				12'd3813	: data1 <= weights[3813];
				12'd3814	: data1 <= weights[3814];
				12'd3815	: data1 <= weights[3815];
				12'd3816	: data1 <= weights[3816];
				12'd3817	: data1 <= weights[3817];
				12'd3818	: data1 <= weights[3818];
				12'd3819	: data1 <= weights[3819];
				12'd3820	: data1 <= weights[3820];
				12'd3821	: data1 <= weights[3821];
				12'd3822	: data1 <= weights[3822];
				12'd3823	: data1 <= weights[3823];
				12'd3824	: data1 <= weights[3824];
				12'd3825	: data1 <= weights[3825];
				12'd3826	: data1 <= weights[3826];
				12'd3827	: data1 <= weights[3827];
				12'd3828	: data1 <= weights[3828];
				12'd3829	: data1 <= weights[3829];
				12'd3830	: data1 <= weights[3830];
				12'd3831	: data1 <= weights[3831];
				12'd3832	: data1 <= weights[3832];
				12'd3833	: data1 <= weights[3833];
				12'd3834	: data1 <= weights[3834];
				12'd3835	: data1 <= weights[3835];
				12'd3836	: data1 <= weights[3836];
				12'd3837	: data1 <= weights[3837];
				12'd3838	: data1 <= weights[3838];
				12'd3839	: data1 <= weights[3839];
				12'd3840	: data1 <= weights[3840];
				12'd3841	: data1 <= weights[3841];
				12'd3842	: data1 <= weights[3842];
				12'd3843	: data1 <= weights[3843];
				12'd3844	: data1 <= weights[3844];
				12'd3845	: data1 <= weights[3845];
				12'd3846	: data1 <= weights[3846];
				12'd3847	: data1 <= weights[3847];
				12'd3848	: data1 <= weights[3848];
				12'd3849	: data1 <= weights[3849];
				12'd3850	: data1 <= weights[3850];
				12'd3851	: data1 <= weights[3851];
				12'd3852	: data1 <= weights[3852];
				12'd3853	: data1 <= weights[3853];
				12'd3854	: data1 <= weights[3854];
				12'd3855	: data1 <= weights[3855];
				12'd3856	: data1 <= weights[3856];
				12'd3857	: data1 <= weights[3857];
				12'd3858	: data1 <= weights[3858];
				12'd3859	: data1 <= weights[3859];
				12'd3860	: data1 <= weights[3860];
				12'd3861	: data1 <= weights[3861];
				12'd3862	: data1 <= weights[3862];
				12'd3863	: data1 <= weights[3863];
				12'd3864	: data1 <= weights[3864];
				12'd3865	: data1 <= weights[3865];
				12'd3866	: data1 <= weights[3866];
				12'd3867	: data1 <= weights[3867];
				12'd3868	: data1 <= weights[3868];
				12'd3869	: data1 <= weights[3869];
				12'd3870	: data1 <= weights[3870];
				12'd3871	: data1 <= weights[3871];
				12'd3872	: data1 <= weights[3872];
				12'd3873	: data1 <= weights[3873];
				12'd3874	: data1 <= weights[3874];
				12'd3875	: data1 <= weights[3875];
				12'd3876	: data1 <= weights[3876];
				12'd3877	: data1 <= weights[3877];
				12'd3878	: data1 <= weights[3878];
				12'd3879	: data1 <= weights[3879];
				12'd3880	: data1 <= weights[3880];
				12'd3881	: data1 <= weights[3881];
				12'd3882	: data1 <= weights[3882];
				12'd3883	: data1 <= weights[3883];
				12'd3884	: data1 <= weights[3884];
				12'd3885	: data1 <= weights[3885];
				12'd3886	: data1 <= weights[3886];
				12'd3887	: data1 <= weights[3887];
				12'd3888	: data1 <= weights[3888];
				12'd3889	: data1 <= weights[3889];
				12'd3890	: data1 <= weights[3890];
				12'd3891	: data1 <= weights[3891];
				12'd3892	: data1 <= weights[3892];
				12'd3893	: data1 <= weights[3893];
				12'd3894	: data1 <= weights[3894];
				12'd3895	: data1 <= weights[3895];
				12'd3896	: data1 <= weights[3896];
				12'd3897	: data1 <= weights[3897];
				12'd3898	: data1 <= weights[3898];
				12'd3899	: data1 <= weights[3899];
				12'd3900	: data1 <= weights[3900];
				12'd3901	: data1 <= weights[3901];
				12'd3902	: data1 <= weights[3902];
				12'd3903	: data1 <= weights[3903];
				12'd3904	: data1 <= weights[3904];
				12'd3905	: data1 <= weights[3905];
				12'd3906	: data1 <= weights[3906];
				12'd3907	: data1 <= weights[3907];
				12'd3908	: data1 <= weights[3908];
				12'd3909	: data1 <= weights[3909];
				12'd3910	: data1 <= weights[3910];
				12'd3911	: data1 <= weights[3911];
				12'd3912	: data1 <= weights[3912];
				12'd3913	: data1 <= weights[3913];
				12'd3914	: data1 <= weights[3914];
				12'd3915	: data1 <= weights[3915];
				12'd3916	: data1 <= weights[3916];
				12'd3917	: data1 <= weights[3917];
				12'd3918	: data1 <= weights[3918];
				12'd3919	: data1 <= weights[3919];
				12'd3920	: data1 <= weights[3920];
				12'd3921	: data1 <= weights[3921];
				12'd3922	: data1 <= weights[3922];
				12'd3923	: data1 <= weights[3923];
				12'd3924	: data1 <= weights[3924];
				12'd3925	: data1 <= weights[3925];
				12'd3926	: data1 <= weights[3926];
				12'd3927	: data1 <= weights[3927];
				12'd3928	: data1 <= weights[3928];
				12'd3929	: data1 <= weights[3929];
				12'd3930	: data1 <= weights[3930];
				12'd3931	: data1 <= weights[3931];
				12'd3932	: data1 <= weights[3932];
				12'd3933	: data1 <= weights[3933];
				12'd3934	: data1 <= weights[3934];
				12'd3935	: data1 <= weights[3935];
				12'd3936	: data1 <= weights[3936];
				12'd3937	: data1 <= weights[3937];
				12'd3938	: data1 <= weights[3938];
				12'd3939	: data1 <= weights[3939];
				12'd3940	: data1 <= weights[3940];
				12'd3941	: data1 <= weights[3941];
				12'd3942	: data1 <= weights[3942];
				12'd3943	: data1 <= weights[3943];
				12'd3944	: data1 <= weights[3944];
				12'd3945	: data1 <= weights[3945];
				12'd3946	: data1 <= weights[3946];
				12'd3947	: data1 <= weights[3947];
				12'd3948	: data1 <= weights[3948];
				12'd3949	: data1 <= weights[3949];
				12'd3950	: data1 <= weights[3950];
				12'd3951	: data1 <= weights[3951];
				12'd3952	: data1 <= weights[3952];
				12'd3953	: data1 <= weights[3953];
				12'd3954	: data1 <= weights[3954];
				12'd3955	: data1 <= weights[3955];
				12'd3956	: data1 <= weights[3956];
				12'd3957	: data1 <= weights[3957];
				12'd3958	: data1 <= weights[3958];
				12'd3959	: data1 <= weights[3959];
				12'd3960	: data1 <= weights[3960];
				12'd3961	: data1 <= weights[3961];
				12'd3962	: data1 <= weights[3962];
				12'd3963	: data1 <= weights[3963];
				12'd3964	: data1 <= weights[3964];
				12'd3965	: data1 <= weights[3965];
				12'd3966	: data1 <= weights[3966];
				12'd3967	: data1 <= weights[3967];
				12'd3968	: data1 <= weights[3968];
				12'd3969	: data1 <= weights[3969];
				12'd3970	: data1 <= weights[3970];
				12'd3971	: data1 <= weights[3971];
				12'd3972	: data1 <= weights[3972];
				12'd3973	: data1 <= weights[3973];
				12'd3974	: data1 <= weights[3974];
				12'd3975	: data1 <= weights[3975];
				12'd3976	: data1 <= weights[3976];
				12'd3977	: data1 <= weights[3977];
				12'd3978	: data1 <= weights[3978];
				12'd3979	: data1 <= weights[3979];
				12'd3980	: data1 <= weights[3980];
				12'd3981	: data1 <= weights[3981];
				12'd3982	: data1 <= weights[3982];
				12'd3983	: data1 <= weights[3983];
				12'd3984	: data1 <= weights[3984];
				12'd3985	: data1 <= weights[3985];
				12'd3986	: data1 <= weights[3986];
				12'd3987	: data1 <= weights[3987];
				12'd3988	: data1 <= weights[3988];
				12'd3989	: data1 <= weights[3989];
				12'd3990	: data1 <= weights[3990];
				12'd3991	: data1 <= weights[3991];
				12'd3992	: data1 <= weights[3992];
				12'd3993	: data1 <= weights[3993];
				12'd3994	: data1 <= weights[3994];
				12'd3995	: data1 <= weights[3995];
				12'd3996	: data1 <= weights[3996];
				12'd3997	: data1 <= weights[3997];
				12'd3998	: data1 <= weights[3998];
				12'd3999	: data1 <= weights[3999];
				12'd4000	: data1 <= weights[4000];
				12'd4001	: data1 <= weights[4001];
				12'd4002	: data1 <= weights[4002];
				12'd4003	: data1 <= weights[4003];
				12'd4004	: data1 <= weights[4004];
				12'd4005	: data1 <= weights[4005];
				12'd4006	: data1 <= weights[4006];
				12'd4007	: data1 <= weights[4007];
				12'd4008	: data1 <= weights[4008];
				12'd4009	: data1 <= weights[4009];
				12'd4010	: data1 <= weights[4010];
				12'd4011	: data1 <= weights[4011];
				12'd4012	: data1 <= weights[4012];
				12'd4013	: data1 <= weights[4013];
				12'd4014	: data1 <= weights[4014];
				12'd4015	: data1 <= weights[4015];
				12'd4016	: data1 <= weights[4016];
				12'd4017	: data1 <= weights[4017];
				12'd4018	: data1 <= weights[4018];
				12'd4019	: data1 <= weights[4019];
				12'd4020	: data1 <= weights[4020];
				12'd4021	: data1 <= weights[4021];
				12'd4022	: data1 <= weights[4022];
				12'd4023	: data1 <= weights[4023];
				12'd4024	: data1 <= weights[4024];
				12'd4025	: data1 <= weights[4025];
				12'd4026	: data1 <= weights[4026];
				12'd4027	: data1 <= weights[4027];
				12'd4028	: data1 <= weights[4028];
				12'd4029	: data1 <= weights[4029];
				12'd4030	: data1 <= weights[4030];
				12'd4031	: data1 <= weights[4031];
				12'd4032	: data1 <= weights[4032];
				12'd4033	: data1 <= weights[4033];
				12'd4034	: data1 <= weights[4034];
				12'd4035	: data1 <= weights[4035];
				12'd4036	: data1 <= weights[4036];
				12'd4037	: data1 <= weights[4037];
				12'd4038	: data1 <= weights[4038];
				12'd4039	: data1 <= weights[4039];
				12'd4040	: data1 <= weights[4040];
				12'd4041	: data1 <= weights[4041];
				12'd4042	: data1 <= weights[4042];
				12'd4043	: data1 <= weights[4043];
				12'd4044	: data1 <= weights[4044];
				12'd4045	: data1 <= weights[4045];
				12'd4046	: data1 <= weights[4046];
				12'd4047	: data1 <= weights[4047];
				12'd4048	: data1 <= weights[4048];
				12'd4049	: data1 <= weights[4049];
				12'd4050	: data1 <= weights[4050];
				default		: data1 <= 16'd0;
			endcase
		end else begin
			data1 <= data1;
		end
	end


	always @(negedge(clk)) begin
		if(enable) begin
			case(address)
				12'd0		: data2 <= weights[1];
				12'd1		: data2 <= weights[2];
				12'd2		: data2 <= weights[3];
				12'd3		: data2 <= weights[4];
				12'd4		: data2 <= weights[5];
				12'd5		: data2 <= weights[6];
				12'd6		: data2 <= weights[7];
				12'd7		: data2 <= weights[8];
				12'd8		: data2 <= weights[9];
				12'd9		: data2 <= weights[10];
				12'd10		: data2 <= weights[11];
				12'd11		: data2 <= weights[12];
				12'd12		: data2 <= weights[13];
				12'd13		: data2 <= weights[14];
				12'd14		: data2 <= weights[15];
				12'd15		: data2 <= weights[16];
				12'd16		: data2 <= weights[17];
				12'd17		: data2 <= weights[18];
				12'd18		: data2 <= weights[19];
				12'd19		: data2 <= weights[20];
				12'd20		: data2 <= weights[21];
				12'd21		: data2 <= weights[22];
				12'd22		: data2 <= weights[23];
				12'd23		: data2 <= weights[24];
				12'd24		: data2 <= weights[25];
				12'd25		: data2 <= weights[26];
				12'd26		: data2 <= weights[27];
				12'd27		: data2 <= weights[28];
				12'd28		: data2 <= weights[29];
				12'd29		: data2 <= weights[30];
				12'd30		: data2 <= weights[31];
				12'd31		: data2 <= weights[32];
				12'd32		: data2 <= weights[33];
				12'd33		: data2 <= weights[34];
				12'd34		: data2 <= weights[35];
				12'd35		: data2 <= weights[36];
				12'd36		: data2 <= weights[37];
				12'd37		: data2 <= weights[38];
				12'd38		: data2 <= weights[39];
				12'd39		: data2 <= weights[40];
				12'd40		: data2 <= weights[41];
				12'd41		: data2 <= weights[42];
				12'd42		: data2 <= weights[43];
				12'd43		: data2 <= weights[44];
				12'd44		: data2 <= weights[45];
				12'd45		: data2 <= weights[46];
				12'd46		: data2 <= weights[47];
				12'd47		: data2 <= weights[48];
				12'd48		: data2 <= weights[49];
				12'd49		: data2 <= weights[50];
				12'd50		: data2 <= weights[51];
				12'd51		: data2 <= weights[52];
				12'd52		: data2 <= weights[53];
				12'd53		: data2 <= weights[54];
				12'd54		: data2 <= weights[55];
				12'd55		: data2 <= weights[56];
				12'd56		: data2 <= weights[57];
				12'd57		: data2 <= weights[58];
				12'd58		: data2 <= weights[59];
				12'd59		: data2 <= weights[60];
				12'd60		: data2 <= weights[61];
				12'd61		: data2 <= weights[62];
				12'd62		: data2 <= weights[63];
				12'd63		: data2 <= weights[64];
				12'd64		: data2 <= weights[65];
				12'd65		: data2 <= weights[66];
				12'd66		: data2 <= weights[67];
				12'd67		: data2 <= weights[68];
				12'd68		: data2 <= weights[69];
				12'd69		: data2 <= weights[70];
				12'd70		: data2 <= weights[71];
				12'd71		: data2 <= weights[72];
				12'd72		: data2 <= weights[73];
				12'd73		: data2 <= weights[74];
				12'd74		: data2 <= weights[75];
				12'd75		: data2 <= weights[76];
				12'd76		: data2 <= weights[77];
				12'd77		: data2 <= weights[78];
				12'd78		: data2 <= weights[79];
				12'd79		: data2 <= weights[80];
				12'd80		: data2 <= weights[81];
				12'd81		: data2 <= weights[82];
				12'd82		: data2 <= weights[83];
				12'd83		: data2 <= weights[84];
				12'd84		: data2 <= weights[85];
				12'd85		: data2 <= weights[86];
				12'd86		: data2 <= weights[87];
				12'd87		: data2 <= weights[88];
				12'd88		: data2 <= weights[89];
				12'd89		: data2 <= weights[90];
				12'd90		: data2 <= weights[91];
				12'd91		: data2 <= weights[92];
				12'd92		: data2 <= weights[93];
				12'd93		: data2 <= weights[94];
				12'd94		: data2 <= weights[95];
				12'd95		: data2 <= weights[96];
				12'd96		: data2 <= weights[97];
				12'd97		: data2 <= weights[98];
				12'd98		: data2 <= weights[99];
				12'd99		: data2 <= weights[100];
				12'd100		: data2 <= weights[101];
				12'd101		: data2 <= weights[102];
				12'd102		: data2 <= weights[103];
				12'd103		: data2 <= weights[104];
				12'd104		: data2 <= weights[105];
				12'd105		: data2 <= weights[106];
				12'd106		: data2 <= weights[107];
				12'd107		: data2 <= weights[108];
				12'd108		: data2 <= weights[109];
				12'd109		: data2 <= weights[110];
				12'd110		: data2 <= weights[111];
				12'd111		: data2 <= weights[112];
				12'd112		: data2 <= weights[113];
				12'd113		: data2 <= weights[114];
				12'd114		: data2 <= weights[115];
				12'd115		: data2 <= weights[116];
				12'd116		: data2 <= weights[117];
				12'd117		: data2 <= weights[118];
				12'd118		: data2 <= weights[119];
				12'd119		: data2 <= weights[120];
				12'd120		: data2 <= weights[121];
				12'd121		: data2 <= weights[122];
				12'd122		: data2 <= weights[123];
				12'd123		: data2 <= weights[124];
				12'd124		: data2 <= weights[125];
				12'd125		: data2 <= weights[126];
				12'd126		: data2 <= weights[127];
				12'd127		: data2 <= weights[128];
				12'd128		: data2 <= weights[129];
				12'd129		: data2 <= weights[130];
				12'd130		: data2 <= weights[131];
				12'd131		: data2 <= weights[132];
				12'd132		: data2 <= weights[133];
				12'd133		: data2 <= weights[134];
				12'd134		: data2 <= weights[135];
				12'd135		: data2 <= weights[136];
				12'd136		: data2 <= weights[137];
				12'd137		: data2 <= weights[138];
				12'd138		: data2 <= weights[139];
				12'd139		: data2 <= weights[140];
				12'd140		: data2 <= weights[141];
				12'd141		: data2 <= weights[142];
				12'd142		: data2 <= weights[143];
				12'd143		: data2 <= weights[144];
				12'd144		: data2 <= weights[145];
				12'd145		: data2 <= weights[146];
				12'd146		: data2 <= weights[147];
				12'd147		: data2 <= weights[148];
				12'd148		: data2 <= weights[149];
				12'd149		: data2 <= weights[150];
				12'd150		: data2 <= weights[151];
				12'd151		: data2 <= weights[152];
				12'd152		: data2 <= weights[153];
				12'd153		: data2 <= weights[154];
				12'd154		: data2 <= weights[155];
				12'd155		: data2 <= weights[156];
				12'd156		: data2 <= weights[157];
				12'd157		: data2 <= weights[158];
				12'd158		: data2 <= weights[159];
				12'd159		: data2 <= weights[160];
				12'd160		: data2 <= weights[161];
				12'd161		: data2 <= weights[162];
				12'd162		: data2 <= weights[163];
				12'd163		: data2 <= weights[164];
				12'd164		: data2 <= weights[165];
				12'd165		: data2 <= weights[166];
				12'd166		: data2 <= weights[167];
				12'd167		: data2 <= weights[168];
				12'd168		: data2 <= weights[169];
				12'd169		: data2 <= weights[170];
				12'd170		: data2 <= weights[171];
				12'd171		: data2 <= weights[172];
				12'd172		: data2 <= weights[173];
				12'd173		: data2 <= weights[174];
				12'd174		: data2 <= weights[175];
				12'd175		: data2 <= weights[176];
				12'd176		: data2 <= weights[177];
				12'd177		: data2 <= weights[178];
				12'd178		: data2 <= weights[179];
				12'd179		: data2 <= weights[180];
				12'd180		: data2 <= weights[181];
				12'd181		: data2 <= weights[182];
				12'd182		: data2 <= weights[183];
				12'd183		: data2 <= weights[184];
				12'd184		: data2 <= weights[185];
				12'd185		: data2 <= weights[186];
				12'd186		: data2 <= weights[187];
				12'd187		: data2 <= weights[188];
				12'd188		: data2 <= weights[189];
				12'd189		: data2 <= weights[190];
				12'd190		: data2 <= weights[191];
				12'd191		: data2 <= weights[192];
				12'd192		: data2 <= weights[193];
				12'd193		: data2 <= weights[194];
				12'd194		: data2 <= weights[195];
				12'd195		: data2 <= weights[196];
				12'd196		: data2 <= weights[197];
				12'd197		: data2 <= weights[198];
				12'd198		: data2 <= weights[199];
				12'd199		: data2 <= weights[200];
				12'd200		: data2 <= weights[201];
				12'd201		: data2 <= weights[202];
				12'd202		: data2 <= weights[203];
				12'd203		: data2 <= weights[204];
				12'd204		: data2 <= weights[205];
				12'd205		: data2 <= weights[206];
				12'd206		: data2 <= weights[207];
				12'd207		: data2 <= weights[208];
				12'd208		: data2 <= weights[209];
				12'd209		: data2 <= weights[210];
				12'd210		: data2 <= weights[211];
				12'd211		: data2 <= weights[212];
				12'd212		: data2 <= weights[213];
				12'd213		: data2 <= weights[214];
				12'd214		: data2 <= weights[215];
				12'd215		: data2 <= weights[216];
				12'd216		: data2 <= weights[217];
				12'd217		: data2 <= weights[218];
				12'd218		: data2 <= weights[219];
				12'd219		: data2 <= weights[220];
				12'd220		: data2 <= weights[221];
				12'd221		: data2 <= weights[222];
				12'd222		: data2 <= weights[223];
				12'd223		: data2 <= weights[224];
				12'd224		: data2 <= weights[225];
				12'd225		: data2 <= weights[226];
				12'd226		: data2 <= weights[227];
				12'd227		: data2 <= weights[228];
				12'd228		: data2 <= weights[229];
				12'd229		: data2 <= weights[230];
				12'd230		: data2 <= weights[231];
				12'd231		: data2 <= weights[232];
				12'd232		: data2 <= weights[233];
				12'd233		: data2 <= weights[234];
				12'd234		: data2 <= weights[235];
				12'd235		: data2 <= weights[236];
				12'd236		: data2 <= weights[237];
				12'd237		: data2 <= weights[238];
				12'd238		: data2 <= weights[239];
				12'd239		: data2 <= weights[240];
				12'd240		: data2 <= weights[241];
				12'd241		: data2 <= weights[242];
				12'd242		: data2 <= weights[243];
				12'd243		: data2 <= weights[244];
				12'd244		: data2 <= weights[245];
				12'd245		: data2 <= weights[246];
				12'd246		: data2 <= weights[247];
				12'd247		: data2 <= weights[248];
				12'd248		: data2 <= weights[249];
				12'd249		: data2 <= weights[250];
				12'd250		: data2 <= weights[251];
				12'd251		: data2 <= weights[252];
				12'd252		: data2 <= weights[253];
				12'd253		: data2 <= weights[254];
				12'd254		: data2 <= weights[255];
				12'd255		: data2 <= weights[256];
				12'd256		: data2 <= weights[257];
				12'd257		: data2 <= weights[258];
				12'd258		: data2 <= weights[259];
				12'd259		: data2 <= weights[260];
				12'd260		: data2 <= weights[261];
				12'd261		: data2 <= weights[262];
				12'd262		: data2 <= weights[263];
				12'd263		: data2 <= weights[264];
				12'd264		: data2 <= weights[265];
				12'd265		: data2 <= weights[266];
				12'd266		: data2 <= weights[267];
				12'd267		: data2 <= weights[268];
				12'd268		: data2 <= weights[269];
				12'd269		: data2 <= weights[270];
				12'd270		: data2 <= weights[271];
				12'd271		: data2 <= weights[272];
				12'd272		: data2 <= weights[273];
				12'd273		: data2 <= weights[274];
				12'd274		: data2 <= weights[275];
				12'd275		: data2 <= weights[276];
				12'd276		: data2 <= weights[277];
				12'd277		: data2 <= weights[278];
				12'd278		: data2 <= weights[279];
				12'd279		: data2 <= weights[280];
				12'd280		: data2 <= weights[281];
				12'd281		: data2 <= weights[282];
				12'd282		: data2 <= weights[283];
				12'd283		: data2 <= weights[284];
				12'd284		: data2 <= weights[285];
				12'd285		: data2 <= weights[286];
				12'd286		: data2 <= weights[287];
				12'd287		: data2 <= weights[288];
				12'd288		: data2 <= weights[289];
				12'd289		: data2 <= weights[290];
				12'd290		: data2 <= weights[291];
				12'd291		: data2 <= weights[292];
				12'd292		: data2 <= weights[293];
				12'd293		: data2 <= weights[294];
				12'd294		: data2 <= weights[295];
				12'd295		: data2 <= weights[296];
				12'd296		: data2 <= weights[297];
				12'd297		: data2 <= weights[298];
				12'd298		: data2 <= weights[299];
				12'd299		: data2 <= weights[300];
				12'd300		: data2 <= weights[301];
				12'd301		: data2 <= weights[302];
				12'd302		: data2 <= weights[303];
				12'd303		: data2 <= weights[304];
				12'd304		: data2 <= weights[305];
				12'd305		: data2 <= weights[306];
				12'd306		: data2 <= weights[307];
				12'd307		: data2 <= weights[308];
				12'd308		: data2 <= weights[309];
				12'd309		: data2 <= weights[310];
				12'd310		: data2 <= weights[311];
				12'd311		: data2 <= weights[312];
				12'd312		: data2 <= weights[313];
				12'd313		: data2 <= weights[314];
				12'd314		: data2 <= weights[315];
				12'd315		: data2 <= weights[316];
				12'd316		: data2 <= weights[317];
				12'd317		: data2 <= weights[318];
				12'd318		: data2 <= weights[319];
				12'd319		: data2 <= weights[320];
				12'd320		: data2 <= weights[321];
				12'd321		: data2 <= weights[322];
				12'd322		: data2 <= weights[323];
				12'd323		: data2 <= weights[324];
				12'd324		: data2 <= weights[325];
				12'd325		: data2 <= weights[326];
				12'd326		: data2 <= weights[327];
				12'd327		: data2 <= weights[328];
				12'd328		: data2 <= weights[329];
				12'd329		: data2 <= weights[330];
				12'd330		: data2 <= weights[331];
				12'd331		: data2 <= weights[332];
				12'd332		: data2 <= weights[333];
				12'd333		: data2 <= weights[334];
				12'd334		: data2 <= weights[335];
				12'd335		: data2 <= weights[336];
				12'd336		: data2 <= weights[337];
				12'd337		: data2 <= weights[338];
				12'd338		: data2 <= weights[339];
				12'd339		: data2 <= weights[340];
				12'd340		: data2 <= weights[341];
				12'd341		: data2 <= weights[342];
				12'd342		: data2 <= weights[343];
				12'd343		: data2 <= weights[344];
				12'd344		: data2 <= weights[345];
				12'd345		: data2 <= weights[346];
				12'd346		: data2 <= weights[347];
				12'd347		: data2 <= weights[348];
				12'd348		: data2 <= weights[349];
				12'd349		: data2 <= weights[350];
				12'd350		: data2 <= weights[351];
				12'd351		: data2 <= weights[352];
				12'd352		: data2 <= weights[353];
				12'd353		: data2 <= weights[354];
				12'd354		: data2 <= weights[355];
				12'd355		: data2 <= weights[356];
				12'd356		: data2 <= weights[357];
				12'd357		: data2 <= weights[358];
				12'd358		: data2 <= weights[359];
				12'd359		: data2 <= weights[360];
				12'd360		: data2 <= weights[361];
				12'd361		: data2 <= weights[362];
				12'd362		: data2 <= weights[363];
				12'd363		: data2 <= weights[364];
				12'd364		: data2 <= weights[365];
				12'd365		: data2 <= weights[366];
				12'd366		: data2 <= weights[367];
				12'd367		: data2 <= weights[368];
				12'd368		: data2 <= weights[369];
				12'd369		: data2 <= weights[370];
				12'd370		: data2 <= weights[371];
				12'd371		: data2 <= weights[372];
				12'd372		: data2 <= weights[373];
				12'd373		: data2 <= weights[374];
				12'd374		: data2 <= weights[375];
				12'd375		: data2 <= weights[376];
				12'd376		: data2 <= weights[377];
				12'd377		: data2 <= weights[378];
				12'd378		: data2 <= weights[379];
				12'd379		: data2 <= weights[380];
				12'd380		: data2 <= weights[381];
				12'd381		: data2 <= weights[382];
				12'd382		: data2 <= weights[383];
				12'd383		: data2 <= weights[384];
				12'd384		: data2 <= weights[385];
				12'd385		: data2 <= weights[386];
				12'd386		: data2 <= weights[387];
				12'd387		: data2 <= weights[388];
				12'd388		: data2 <= weights[389];
				12'd389		: data2 <= weights[390];
				12'd390		: data2 <= weights[391];
				12'd391		: data2 <= weights[392];
				12'd392		: data2 <= weights[393];
				12'd393		: data2 <= weights[394];
				12'd394		: data2 <= weights[395];
				12'd395		: data2 <= weights[396];
				12'd396		: data2 <= weights[397];
				12'd397		: data2 <= weights[398];
				12'd398		: data2 <= weights[399];
				12'd399		: data2 <= weights[400];
				12'd400		: data2 <= weights[401];
				12'd401		: data2 <= weights[402];
				12'd402		: data2 <= weights[403];
				12'd403		: data2 <= weights[404];
				12'd404		: data2 <= weights[405];
				12'd405		: data2 <= weights[406];
				12'd406		: data2 <= weights[407];
				12'd407		: data2 <= weights[408];
				12'd408		: data2 <= weights[409];
				12'd409		: data2 <= weights[410];
				12'd410		: data2 <= weights[411];
				12'd411		: data2 <= weights[412];
				12'd412		: data2 <= weights[413];
				12'd413		: data2 <= weights[414];
				12'd414		: data2 <= weights[415];
				12'd415		: data2 <= weights[416];
				12'd416		: data2 <= weights[417];
				12'd417		: data2 <= weights[418];
				12'd418		: data2 <= weights[419];
				12'd419		: data2 <= weights[420];
				12'd420		: data2 <= weights[421];
				12'd421		: data2 <= weights[422];
				12'd422		: data2 <= weights[423];
				12'd423		: data2 <= weights[424];
				12'd424		: data2 <= weights[425];
				12'd425		: data2 <= weights[426];
				12'd426		: data2 <= weights[427];
				12'd427		: data2 <= weights[428];
				12'd428		: data2 <= weights[429];
				12'd429		: data2 <= weights[430];
				12'd430		: data2 <= weights[431];
				12'd431		: data2 <= weights[432];
				12'd432		: data2 <= weights[433];
				12'd433		: data2 <= weights[434];
				12'd434		: data2 <= weights[435];
				12'd435		: data2 <= weights[436];
				12'd436		: data2 <= weights[437];
				12'd437		: data2 <= weights[438];
				12'd438		: data2 <= weights[439];
				12'd439		: data2 <= weights[440];
				12'd440		: data2 <= weights[441];
				12'd441		: data2 <= weights[442];
				12'd442		: data2 <= weights[443];
				12'd443		: data2 <= weights[444];
				12'd444		: data2 <= weights[445];
				12'd445		: data2 <= weights[446];
				12'd446		: data2 <= weights[447];
				12'd447		: data2 <= weights[448];
				12'd448		: data2 <= weights[449];
				12'd449		: data2 <= weights[450];
				12'd450		: data2 <= weights[451];
				12'd451		: data2 <= weights[452];
				12'd452		: data2 <= weights[453];
				12'd453		: data2 <= weights[454];
				12'd454		: data2 <= weights[455];
				12'd455		: data2 <= weights[456];
				12'd456		: data2 <= weights[457];
				12'd457		: data2 <= weights[458];
				12'd458		: data2 <= weights[459];
				12'd459		: data2 <= weights[460];
				12'd460		: data2 <= weights[461];
				12'd461		: data2 <= weights[462];
				12'd462		: data2 <= weights[463];
				12'd463		: data2 <= weights[464];
				12'd464		: data2 <= weights[465];
				12'd465		: data2 <= weights[466];
				12'd466		: data2 <= weights[467];
				12'd467		: data2 <= weights[468];
				12'd468		: data2 <= weights[469];
				12'd469		: data2 <= weights[470];
				12'd470		: data2 <= weights[471];
				12'd471		: data2 <= weights[472];
				12'd472		: data2 <= weights[473];
				12'd473		: data2 <= weights[474];
				12'd474		: data2 <= weights[475];
				12'd475		: data2 <= weights[476];
				12'd476		: data2 <= weights[477];
				12'd477		: data2 <= weights[478];
				12'd478		: data2 <= weights[479];
				12'd479		: data2 <= weights[480];
				12'd480		: data2 <= weights[481];
				12'd481		: data2 <= weights[482];
				12'd482		: data2 <= weights[483];
				12'd483		: data2 <= weights[484];
				12'd484		: data2 <= weights[485];
				12'd485		: data2 <= weights[486];
				12'd486		: data2 <= weights[487];
				12'd487		: data2 <= weights[488];
				12'd488		: data2 <= weights[489];
				12'd489		: data2 <= weights[490];
				12'd490		: data2 <= weights[491];
				12'd491		: data2 <= weights[492];
				12'd492		: data2 <= weights[493];
				12'd493		: data2 <= weights[494];
				12'd494		: data2 <= weights[495];
				12'd495		: data2 <= weights[496];
				12'd496		: data2 <= weights[497];
				12'd497		: data2 <= weights[498];
				12'd498		: data2 <= weights[499];
				12'd499		: data2 <= weights[500];
				12'd500		: data2 <= weights[501];
				12'd501		: data2 <= weights[502];
				12'd502		: data2 <= weights[503];
				12'd503		: data2 <= weights[504];
				12'd504		: data2 <= weights[505];
				12'd505		: data2 <= weights[506];
				12'd506		: data2 <= weights[507];
				12'd507		: data2 <= weights[508];
				12'd508		: data2 <= weights[509];
				12'd509		: data2 <= weights[510];
				12'd510		: data2 <= weights[511];
				12'd511		: data2 <= weights[512];
				12'd512		: data2 <= weights[513];
				12'd513		: data2 <= weights[514];
				12'd514		: data2 <= weights[515];
				12'd515		: data2 <= weights[516];
				12'd516		: data2 <= weights[517];
				12'd517		: data2 <= weights[518];
				12'd518		: data2 <= weights[519];
				12'd519		: data2 <= weights[520];
				12'd520		: data2 <= weights[521];
				12'd521		: data2 <= weights[522];
				12'd522		: data2 <= weights[523];
				12'd523		: data2 <= weights[524];
				12'd524		: data2 <= weights[525];
				12'd525		: data2 <= weights[526];
				12'd526		: data2 <= weights[527];
				12'd527		: data2 <= weights[528];
				12'd528		: data2 <= weights[529];
				12'd529		: data2 <= weights[530];
				12'd530		: data2 <= weights[531];
				12'd531		: data2 <= weights[532];
				12'd532		: data2 <= weights[533];
				12'd533		: data2 <= weights[534];
				12'd534		: data2 <= weights[535];
				12'd535		: data2 <= weights[536];
				12'd536		: data2 <= weights[537];
				12'd537		: data2 <= weights[538];
				12'd538		: data2 <= weights[539];
				12'd539		: data2 <= weights[540];
				12'd540		: data2 <= weights[541];
				12'd541		: data2 <= weights[542];
				12'd542		: data2 <= weights[543];
				12'd543		: data2 <= weights[544];
				12'd544		: data2 <= weights[545];
				12'd545		: data2 <= weights[546];
				12'd546		: data2 <= weights[547];
				12'd547		: data2 <= weights[548];
				12'd548		: data2 <= weights[549];
				12'd549		: data2 <= weights[550];
				12'd550		: data2 <= weights[551];
				12'd551		: data2 <= weights[552];
				12'd552		: data2 <= weights[553];
				12'd553		: data2 <= weights[554];
				12'd554		: data2 <= weights[555];
				12'd555		: data2 <= weights[556];
				12'd556		: data2 <= weights[557];
				12'd557		: data2 <= weights[558];
				12'd558		: data2 <= weights[559];
				12'd559		: data2 <= weights[560];
				12'd560		: data2 <= weights[561];
				12'd561		: data2 <= weights[562];
				12'd562		: data2 <= weights[563];
				12'd563		: data2 <= weights[564];
				12'd564		: data2 <= weights[565];
				12'd565		: data2 <= weights[566];
				12'd566		: data2 <= weights[567];
				12'd567		: data2 <= weights[568];
				12'd568		: data2 <= weights[569];
				12'd569		: data2 <= weights[570];
				12'd570		: data2 <= weights[571];
				12'd571		: data2 <= weights[572];
				12'd572		: data2 <= weights[573];
				12'd573		: data2 <= weights[574];
				12'd574		: data2 <= weights[575];
				12'd575		: data2 <= weights[576];
				12'd576		: data2 <= weights[577];
				12'd577		: data2 <= weights[578];
				12'd578		: data2 <= weights[579];
				12'd579		: data2 <= weights[580];
				12'd580		: data2 <= weights[581];
				12'd581		: data2 <= weights[582];
				12'd582		: data2 <= weights[583];
				12'd583		: data2 <= weights[584];
				12'd584		: data2 <= weights[585];
				12'd585		: data2 <= weights[586];
				12'd586		: data2 <= weights[587];
				12'd587		: data2 <= weights[588];
				12'd588		: data2 <= weights[589];
				12'd589		: data2 <= weights[590];
				12'd590		: data2 <= weights[591];
				12'd591		: data2 <= weights[592];
				12'd592		: data2 <= weights[593];
				12'd593		: data2 <= weights[594];
				12'd594		: data2 <= weights[595];
				12'd595		: data2 <= weights[596];
				12'd596		: data2 <= weights[597];
				12'd597		: data2 <= weights[598];
				12'd598		: data2 <= weights[599];
				12'd599		: data2 <= weights[600];
				12'd600		: data2 <= weights[601];
				12'd601		: data2 <= weights[602];
				12'd602		: data2 <= weights[603];
				12'd603		: data2 <= weights[604];
				12'd604		: data2 <= weights[605];
				12'd605		: data2 <= weights[606];
				12'd606		: data2 <= weights[607];
				12'd607		: data2 <= weights[608];
				12'd608		: data2 <= weights[609];
				12'd609		: data2 <= weights[610];
				12'd610		: data2 <= weights[611];
				12'd611		: data2 <= weights[612];
				12'd612		: data2 <= weights[613];
				12'd613		: data2 <= weights[614];
				12'd614		: data2 <= weights[615];
				12'd615		: data2 <= weights[616];
				12'd616		: data2 <= weights[617];
				12'd617		: data2 <= weights[618];
				12'd618		: data2 <= weights[619];
				12'd619		: data2 <= weights[620];
				12'd620		: data2 <= weights[621];
				12'd621		: data2 <= weights[622];
				12'd622		: data2 <= weights[623];
				12'd623		: data2 <= weights[624];
				12'd624		: data2 <= weights[625];
				12'd625		: data2 <= weights[626];
				12'd626		: data2 <= weights[627];
				12'd627		: data2 <= weights[628];
				12'd628		: data2 <= weights[629];
				12'd629		: data2 <= weights[630];
				12'd630		: data2 <= weights[631];
				12'd631		: data2 <= weights[632];
				12'd632		: data2 <= weights[633];
				12'd633		: data2 <= weights[634];
				12'd634		: data2 <= weights[635];
				12'd635		: data2 <= weights[636];
				12'd636		: data2 <= weights[637];
				12'd637		: data2 <= weights[638];
				12'd638		: data2 <= weights[639];
				12'd639		: data2 <= weights[640];
				12'd640		: data2 <= weights[641];
				12'd641		: data2 <= weights[642];
				12'd642		: data2 <= weights[643];
				12'd643		: data2 <= weights[644];
				12'd644		: data2 <= weights[645];
				12'd645		: data2 <= weights[646];
				12'd646		: data2 <= weights[647];
				12'd647		: data2 <= weights[648];
				12'd648		: data2 <= weights[649];
				12'd649		: data2 <= weights[650];
				12'd650		: data2 <= weights[651];
				12'd651		: data2 <= weights[652];
				12'd652		: data2 <= weights[653];
				12'd653		: data2 <= weights[654];
				12'd654		: data2 <= weights[655];
				12'd655		: data2 <= weights[656];
				12'd656		: data2 <= weights[657];
				12'd657		: data2 <= weights[658];
				12'd658		: data2 <= weights[659];
				12'd659		: data2 <= weights[660];
				12'd660		: data2 <= weights[661];
				12'd661		: data2 <= weights[662];
				12'd662		: data2 <= weights[663];
				12'd663		: data2 <= weights[664];
				12'd664		: data2 <= weights[665];
				12'd665		: data2 <= weights[666];
				12'd666		: data2 <= weights[667];
				12'd667		: data2 <= weights[668];
				12'd668		: data2 <= weights[669];
				12'd669		: data2 <= weights[670];
				12'd670		: data2 <= weights[671];
				12'd671		: data2 <= weights[672];
				12'd672		: data2 <= weights[673];
				12'd673		: data2 <= weights[674];
				12'd674		: data2 <= weights[675];
				12'd675		: data2 <= weights[676];
				12'd676		: data2 <= weights[677];
				12'd677		: data2 <= weights[678];
				12'd678		: data2 <= weights[679];
				12'd679		: data2 <= weights[680];
				12'd680		: data2 <= weights[681];
				12'd681		: data2 <= weights[682];
				12'd682		: data2 <= weights[683];
				12'd683		: data2 <= weights[684];
				12'd684		: data2 <= weights[685];
				12'd685		: data2 <= weights[686];
				12'd686		: data2 <= weights[687];
				12'd687		: data2 <= weights[688];
				12'd688		: data2 <= weights[689];
				12'd689		: data2 <= weights[690];
				12'd690		: data2 <= weights[691];
				12'd691		: data2 <= weights[692];
				12'd692		: data2 <= weights[693];
				12'd693		: data2 <= weights[694];
				12'd694		: data2 <= weights[695];
				12'd695		: data2 <= weights[696];
				12'd696		: data2 <= weights[697];
				12'd697		: data2 <= weights[698];
				12'd698		: data2 <= weights[699];
				12'd699		: data2 <= weights[700];
				12'd700		: data2 <= weights[701];
				12'd701		: data2 <= weights[702];
				12'd702		: data2 <= weights[703];
				12'd703		: data2 <= weights[704];
				12'd704		: data2 <= weights[705];
				12'd705		: data2 <= weights[706];
				12'd706		: data2 <= weights[707];
				12'd707		: data2 <= weights[708];
				12'd708		: data2 <= weights[709];
				12'd709		: data2 <= weights[710];
				12'd710		: data2 <= weights[711];
				12'd711		: data2 <= weights[712];
				12'd712		: data2 <= weights[713];
				12'd713		: data2 <= weights[714];
				12'd714		: data2 <= weights[715];
				12'd715		: data2 <= weights[716];
				12'd716		: data2 <= weights[717];
				12'd717		: data2 <= weights[718];
				12'd718		: data2 <= weights[719];
				12'd719		: data2 <= weights[720];
				12'd720		: data2 <= weights[721];
				12'd721		: data2 <= weights[722];
				12'd722		: data2 <= weights[723];
				12'd723		: data2 <= weights[724];
				12'd724		: data2 <= weights[725];
				12'd725		: data2 <= weights[726];
				12'd726		: data2 <= weights[727];
				12'd727		: data2 <= weights[728];
				12'd728		: data2 <= weights[729];
				12'd729		: data2 <= weights[730];
				12'd730		: data2 <= weights[731];
				12'd731		: data2 <= weights[732];
				12'd732		: data2 <= weights[733];
				12'd733		: data2 <= weights[734];
				12'd734		: data2 <= weights[735];
				12'd735		: data2 <= weights[736];
				12'd736		: data2 <= weights[737];
				12'd737		: data2 <= weights[738];
				12'd738		: data2 <= weights[739];
				12'd739		: data2 <= weights[740];
				12'd740		: data2 <= weights[741];
				12'd741		: data2 <= weights[742];
				12'd742		: data2 <= weights[743];
				12'd743		: data2 <= weights[744];
				12'd744		: data2 <= weights[745];
				12'd745		: data2 <= weights[746];
				12'd746		: data2 <= weights[747];
				12'd747		: data2 <= weights[748];
				12'd748		: data2 <= weights[749];
				12'd749		: data2 <= weights[750];
				12'd750		: data2 <= weights[751];
				12'd751		: data2 <= weights[752];
				12'd752		: data2 <= weights[753];
				12'd753		: data2 <= weights[754];
				12'd754		: data2 <= weights[755];
				12'd755		: data2 <= weights[756];
				12'd756		: data2 <= weights[757];
				12'd757		: data2 <= weights[758];
				12'd758		: data2 <= weights[759];
				12'd759		: data2 <= weights[760];
				12'd760		: data2 <= weights[761];
				12'd761		: data2 <= weights[762];
				12'd762		: data2 <= weights[763];
				12'd763		: data2 <= weights[764];
				12'd764		: data2 <= weights[765];
				12'd765		: data2 <= weights[766];
				12'd766		: data2 <= weights[767];
				12'd767		: data2 <= weights[768];
				12'd768		: data2 <= weights[769];
				12'd769		: data2 <= weights[770];
				12'd770		: data2 <= weights[771];
				12'd771		: data2 <= weights[772];
				12'd772		: data2 <= weights[773];
				12'd773		: data2 <= weights[774];
				12'd774		: data2 <= weights[775];
				12'd775		: data2 <= weights[776];
				12'd776		: data2 <= weights[777];
				12'd777		: data2 <= weights[778];
				12'd778		: data2 <= weights[779];
				12'd779		: data2 <= weights[780];
				12'd780		: data2 <= weights[781];
				12'd781		: data2 <= weights[782];
				12'd782		: data2 <= weights[783];
				12'd783		: data2 <= weights[784];
				12'd784		: data2 <= weights[785];
				12'd785		: data2 <= weights[786];
				12'd786		: data2 <= weights[787];
				12'd787		: data2 <= weights[788];
				12'd788		: data2 <= weights[789];
				12'd789		: data2 <= weights[790];
				12'd790		: data2 <= weights[791];
				12'd791		: data2 <= weights[792];
				12'd792		: data2 <= weights[793];
				12'd793		: data2 <= weights[794];
				12'd794		: data2 <= weights[795];
				12'd795		: data2 <= weights[796];
				12'd796		: data2 <= weights[797];
				12'd797		: data2 <= weights[798];
				12'd798		: data2 <= weights[799];
				12'd799		: data2 <= weights[800];
				12'd800		: data2 <= weights[801];
				12'd801		: data2 <= weights[802];
				12'd802		: data2 <= weights[803];
				12'd803		: data2 <= weights[804];
				12'd804		: data2 <= weights[805];
				12'd805		: data2 <= weights[806];
				12'd806		: data2 <= weights[807];
				12'd807		: data2 <= weights[808];
				12'd808		: data2 <= weights[809];
				12'd809		: data2 <= weights[810];
				12'd810		: data2 <= weights[811];
				12'd811		: data2 <= weights[812];
				12'd812		: data2 <= weights[813];
				12'd813		: data2 <= weights[814];
				12'd814		: data2 <= weights[815];
				12'd815		: data2 <= weights[816];
				12'd816		: data2 <= weights[817];
				12'd817		: data2 <= weights[818];
				12'd818		: data2 <= weights[819];
				12'd819		: data2 <= weights[820];
				12'd820		: data2 <= weights[821];
				12'd821		: data2 <= weights[822];
				12'd822		: data2 <= weights[823];
				12'd823		: data2 <= weights[824];
				12'd824		: data2 <= weights[825];
				12'd825		: data2 <= weights[826];
				12'd826		: data2 <= weights[827];
				12'd827		: data2 <= weights[828];
				12'd828		: data2 <= weights[829];
				12'd829		: data2 <= weights[830];
				12'd830		: data2 <= weights[831];
				12'd831		: data2 <= weights[832];
				12'd832		: data2 <= weights[833];
				12'd833		: data2 <= weights[834];
				12'd834		: data2 <= weights[835];
				12'd835		: data2 <= weights[836];
				12'd836		: data2 <= weights[837];
				12'd837		: data2 <= weights[838];
				12'd838		: data2 <= weights[839];
				12'd839		: data2 <= weights[840];
				12'd840		: data2 <= weights[841];
				12'd841		: data2 <= weights[842];
				12'd842		: data2 <= weights[843];
				12'd843		: data2 <= weights[844];
				12'd844		: data2 <= weights[845];
				12'd845		: data2 <= weights[846];
				12'd846		: data2 <= weights[847];
				12'd847		: data2 <= weights[848];
				12'd848		: data2 <= weights[849];
				12'd849		: data2 <= weights[850];
				12'd850		: data2 <= weights[851];
				12'd851		: data2 <= weights[852];
				12'd852		: data2 <= weights[853];
				12'd853		: data2 <= weights[854];
				12'd854		: data2 <= weights[855];
				12'd855		: data2 <= weights[856];
				12'd856		: data2 <= weights[857];
				12'd857		: data2 <= weights[858];
				12'd858		: data2 <= weights[859];
				12'd859		: data2 <= weights[860];
				12'd860		: data2 <= weights[861];
				12'd861		: data2 <= weights[862];
				12'd862		: data2 <= weights[863];
				12'd863		: data2 <= weights[864];
				12'd864		: data2 <= weights[865];
				12'd865		: data2 <= weights[866];
				12'd866		: data2 <= weights[867];
				12'd867		: data2 <= weights[868];
				12'd868		: data2 <= weights[869];
				12'd869		: data2 <= weights[870];
				12'd870		: data2 <= weights[871];
				12'd871		: data2 <= weights[872];
				12'd872		: data2 <= weights[873];
				12'd873		: data2 <= weights[874];
				12'd874		: data2 <= weights[875];
				12'd875		: data2 <= weights[876];
				12'd876		: data2 <= weights[877];
				12'd877		: data2 <= weights[878];
				12'd878		: data2 <= weights[879];
				12'd879		: data2 <= weights[880];
				12'd880		: data2 <= weights[881];
				12'd881		: data2 <= weights[882];
				12'd882		: data2 <= weights[883];
				12'd883		: data2 <= weights[884];
				12'd884		: data2 <= weights[885];
				12'd885		: data2 <= weights[886];
				12'd886		: data2 <= weights[887];
				12'd887		: data2 <= weights[888];
				12'd888		: data2 <= weights[889];
				12'd889		: data2 <= weights[890];
				12'd890		: data2 <= weights[891];
				12'd891		: data2 <= weights[892];
				12'd892		: data2 <= weights[893];
				12'd893		: data2 <= weights[894];
				12'd894		: data2 <= weights[895];
				12'd895		: data2 <= weights[896];
				12'd896		: data2 <= weights[897];
				12'd897		: data2 <= weights[898];
				12'd898		: data2 <= weights[899];
				12'd899		: data2 <= weights[900];
				12'd900		: data2 <= weights[901];
				12'd901		: data2 <= weights[902];
				12'd902		: data2 <= weights[903];
				12'd903		: data2 <= weights[904];
				12'd904		: data2 <= weights[905];
				12'd905		: data2 <= weights[906];
				12'd906		: data2 <= weights[907];
				12'd907		: data2 <= weights[908];
				12'd908		: data2 <= weights[909];
				12'd909		: data2 <= weights[910];
				12'd910		: data2 <= weights[911];
				12'd911		: data2 <= weights[912];
				12'd912		: data2 <= weights[913];
				12'd913		: data2 <= weights[914];
				12'd914		: data2 <= weights[915];
				12'd915		: data2 <= weights[916];
				12'd916		: data2 <= weights[917];
				12'd917		: data2 <= weights[918];
				12'd918		: data2 <= weights[919];
				12'd919		: data2 <= weights[920];
				12'd920		: data2 <= weights[921];
				12'd921		: data2 <= weights[922];
				12'd922		: data2 <= weights[923];
				12'd923		: data2 <= weights[924];
				12'd924		: data2 <= weights[925];
				12'd925		: data2 <= weights[926];
				12'd926		: data2 <= weights[927];
				12'd927		: data2 <= weights[928];
				12'd928		: data2 <= weights[929];
				12'd929		: data2 <= weights[930];
				12'd930		: data2 <= weights[931];
				12'd931		: data2 <= weights[932];
				12'd932		: data2 <= weights[933];
				12'd933		: data2 <= weights[934];
				12'd934		: data2 <= weights[935];
				12'd935		: data2 <= weights[936];
				12'd936		: data2 <= weights[937];
				12'd937		: data2 <= weights[938];
				12'd938		: data2 <= weights[939];
				12'd939		: data2 <= weights[940];
				12'd940		: data2 <= weights[941];
				12'd941		: data2 <= weights[942];
				12'd942		: data2 <= weights[943];
				12'd943		: data2 <= weights[944];
				12'd944		: data2 <= weights[945];
				12'd945		: data2 <= weights[946];
				12'd946		: data2 <= weights[947];
				12'd947		: data2 <= weights[948];
				12'd948		: data2 <= weights[949];
				12'd949		: data2 <= weights[950];
				12'd950		: data2 <= weights[951];
				12'd951		: data2 <= weights[952];
				12'd952		: data2 <= weights[953];
				12'd953		: data2 <= weights[954];
				12'd954		: data2 <= weights[955];
				12'd955		: data2 <= weights[956];
				12'd956		: data2 <= weights[957];
				12'd957		: data2 <= weights[958];
				12'd958		: data2 <= weights[959];
				12'd959		: data2 <= weights[960];
				12'd960		: data2 <= weights[961];
				12'd961		: data2 <= weights[962];
				12'd962		: data2 <= weights[963];
				12'd963		: data2 <= weights[964];
				12'd964		: data2 <= weights[965];
				12'd965		: data2 <= weights[966];
				12'd966		: data2 <= weights[967];
				12'd967		: data2 <= weights[968];
				12'd968		: data2 <= weights[969];
				12'd969		: data2 <= weights[970];
				12'd970		: data2 <= weights[971];
				12'd971		: data2 <= weights[972];
				12'd972		: data2 <= weights[973];
				12'd973		: data2 <= weights[974];
				12'd974		: data2 <= weights[975];
				12'd975		: data2 <= weights[976];
				12'd976		: data2 <= weights[977];
				12'd977		: data2 <= weights[978];
				12'd978		: data2 <= weights[979];
				12'd979		: data2 <= weights[980];
				12'd980		: data2 <= weights[981];
				12'd981		: data2 <= weights[982];
				12'd982		: data2 <= weights[983];
				12'd983		: data2 <= weights[984];
				12'd984		: data2 <= weights[985];
				12'd985		: data2 <= weights[986];
				12'd986		: data2 <= weights[987];
				12'd987		: data2 <= weights[988];
				12'd988		: data2 <= weights[989];
				12'd989		: data2 <= weights[990];
				12'd990		: data2 <= weights[991];
				12'd991		: data2 <= weights[992];
				12'd992		: data2 <= weights[993];
				12'd993		: data2 <= weights[994];
				12'd994		: data2 <= weights[995];
				12'd995		: data2 <= weights[996];
				12'd996		: data2 <= weights[997];
				12'd997		: data2 <= weights[998];
				12'd998		: data2 <= weights[999];
				12'd999		: data2 <= weights[1000];
				12'd1000	: data2 <= weights[1001];
				12'd1001	: data2 <= weights[1002];
				12'd1002	: data2 <= weights[1003];
				12'd1003	: data2 <= weights[1004];
				12'd1004	: data2 <= weights[1005];
				12'd1005	: data2 <= weights[1006];
				12'd1006	: data2 <= weights[1007];
				12'd1007	: data2 <= weights[1008];
				12'd1008	: data2 <= weights[1009];
				12'd1009	: data2 <= weights[1010];
				12'd1010	: data2 <= weights[1011];
				12'd1011	: data2 <= weights[1012];
				12'd1012	: data2 <= weights[1013];
				12'd1013	: data2 <= weights[1014];
				12'd1014	: data2 <= weights[1015];
				12'd1015	: data2 <= weights[1016];
				12'd1016	: data2 <= weights[1017];
				12'd1017	: data2 <= weights[1018];
				12'd1018	: data2 <= weights[1019];
				12'd1019	: data2 <= weights[1020];
				12'd1020	: data2 <= weights[1021];
				12'd1021	: data2 <= weights[1022];
				12'd1022	: data2 <= weights[1023];
				12'd1023	: data2 <= weights[1024];
				12'd1024	: data2 <= weights[1025];
				12'd1025	: data2 <= weights[1026];
				12'd1026	: data2 <= weights[1027];
				12'd1027	: data2 <= weights[1028];
				12'd1028	: data2 <= weights[1029];
				12'd1029	: data2 <= weights[1030];
				12'd1030	: data2 <= weights[1031];
				12'd1031	: data2 <= weights[1032];
				12'd1032	: data2 <= weights[1033];
				12'd1033	: data2 <= weights[1034];
				12'd1034	: data2 <= weights[1035];
				12'd1035	: data2 <= weights[1036];
				12'd1036	: data2 <= weights[1037];
				12'd1037	: data2 <= weights[1038];
				12'd1038	: data2 <= weights[1039];
				12'd1039	: data2 <= weights[1040];
				12'd1040	: data2 <= weights[1041];
				12'd1041	: data2 <= weights[1042];
				12'd1042	: data2 <= weights[1043];
				12'd1043	: data2 <= weights[1044];
				12'd1044	: data2 <= weights[1045];
				12'd1045	: data2 <= weights[1046];
				12'd1046	: data2 <= weights[1047];
				12'd1047	: data2 <= weights[1048];
				12'd1048	: data2 <= weights[1049];
				12'd1049	: data2 <= weights[1050];
				12'd1050	: data2 <= weights[1051];
				12'd1051	: data2 <= weights[1052];
				12'd1052	: data2 <= weights[1053];
				12'd1053	: data2 <= weights[1054];
				12'd1054	: data2 <= weights[1055];
				12'd1055	: data2 <= weights[1056];
				12'd1056	: data2 <= weights[1057];
				12'd1057	: data2 <= weights[1058];
				12'd1058	: data2 <= weights[1059];
				12'd1059	: data2 <= weights[1060];
				12'd1060	: data2 <= weights[1061];
				12'd1061	: data2 <= weights[1062];
				12'd1062	: data2 <= weights[1063];
				12'd1063	: data2 <= weights[1064];
				12'd1064	: data2 <= weights[1065];
				12'd1065	: data2 <= weights[1066];
				12'd1066	: data2 <= weights[1067];
				12'd1067	: data2 <= weights[1068];
				12'd1068	: data2 <= weights[1069];
				12'd1069	: data2 <= weights[1070];
				12'd1070	: data2 <= weights[1071];
				12'd1071	: data2 <= weights[1072];
				12'd1072	: data2 <= weights[1073];
				12'd1073	: data2 <= weights[1074];
				12'd1074	: data2 <= weights[1075];
				12'd1075	: data2 <= weights[1076];
				12'd1076	: data2 <= weights[1077];
				12'd1077	: data2 <= weights[1078];
				12'd1078	: data2 <= weights[1079];
				12'd1079	: data2 <= weights[1080];
				12'd1080	: data2 <= weights[1081];
				12'd1081	: data2 <= weights[1082];
				12'd1082	: data2 <= weights[1083];
				12'd1083	: data2 <= weights[1084];
				12'd1084	: data2 <= weights[1085];
				12'd1085	: data2 <= weights[1086];
				12'd1086	: data2 <= weights[1087];
				12'd1087	: data2 <= weights[1088];
				12'd1088	: data2 <= weights[1089];
				12'd1089	: data2 <= weights[1090];
				12'd1090	: data2 <= weights[1091];
				12'd1091	: data2 <= weights[1092];
				12'd1092	: data2 <= weights[1093];
				12'd1093	: data2 <= weights[1094];
				12'd1094	: data2 <= weights[1095];
				12'd1095	: data2 <= weights[1096];
				12'd1096	: data2 <= weights[1097];
				12'd1097	: data2 <= weights[1098];
				12'd1098	: data2 <= weights[1099];
				12'd1099	: data2 <= weights[1100];
				12'd1100	: data2 <= weights[1101];
				12'd1101	: data2 <= weights[1102];
				12'd1102	: data2 <= weights[1103];
				12'd1103	: data2 <= weights[1104];
				12'd1104	: data2 <= weights[1105];
				12'd1105	: data2 <= weights[1106];
				12'd1106	: data2 <= weights[1107];
				12'd1107	: data2 <= weights[1108];
				12'd1108	: data2 <= weights[1109];
				12'd1109	: data2 <= weights[1110];
				12'd1110	: data2 <= weights[1111];
				12'd1111	: data2 <= weights[1112];
				12'd1112	: data2 <= weights[1113];
				12'd1113	: data2 <= weights[1114];
				12'd1114	: data2 <= weights[1115];
				12'd1115	: data2 <= weights[1116];
				12'd1116	: data2 <= weights[1117];
				12'd1117	: data2 <= weights[1118];
				12'd1118	: data2 <= weights[1119];
				12'd1119	: data2 <= weights[1120];
				12'd1120	: data2 <= weights[1121];
				12'd1121	: data2 <= weights[1122];
				12'd1122	: data2 <= weights[1123];
				12'd1123	: data2 <= weights[1124];
				12'd1124	: data2 <= weights[1125];
				12'd1125	: data2 <= weights[1126];
				12'd1126	: data2 <= weights[1127];
				12'd1127	: data2 <= weights[1128];
				12'd1128	: data2 <= weights[1129];
				12'd1129	: data2 <= weights[1130];
				12'd1130	: data2 <= weights[1131];
				12'd1131	: data2 <= weights[1132];
				12'd1132	: data2 <= weights[1133];
				12'd1133	: data2 <= weights[1134];
				12'd1134	: data2 <= weights[1135];
				12'd1135	: data2 <= weights[1136];
				12'd1136	: data2 <= weights[1137];
				12'd1137	: data2 <= weights[1138];
				12'd1138	: data2 <= weights[1139];
				12'd1139	: data2 <= weights[1140];
				12'd1140	: data2 <= weights[1141];
				12'd1141	: data2 <= weights[1142];
				12'd1142	: data2 <= weights[1143];
				12'd1143	: data2 <= weights[1144];
				12'd1144	: data2 <= weights[1145];
				12'd1145	: data2 <= weights[1146];
				12'd1146	: data2 <= weights[1147];
				12'd1147	: data2 <= weights[1148];
				12'd1148	: data2 <= weights[1149];
				12'd1149	: data2 <= weights[1150];
				12'd1150	: data2 <= weights[1151];
				12'd1151	: data2 <= weights[1152];
				12'd1152	: data2 <= weights[1153];
				12'd1153	: data2 <= weights[1154];
				12'd1154	: data2 <= weights[1155];
				12'd1155	: data2 <= weights[1156];
				12'd1156	: data2 <= weights[1157];
				12'd1157	: data2 <= weights[1158];
				12'd1158	: data2 <= weights[1159];
				12'd1159	: data2 <= weights[1160];
				12'd1160	: data2 <= weights[1161];
				12'd1161	: data2 <= weights[1162];
				12'd1162	: data2 <= weights[1163];
				12'd1163	: data2 <= weights[1164];
				12'd1164	: data2 <= weights[1165];
				12'd1165	: data2 <= weights[1166];
				12'd1166	: data2 <= weights[1167];
				12'd1167	: data2 <= weights[1168];
				12'd1168	: data2 <= weights[1169];
				12'd1169	: data2 <= weights[1170];
				12'd1170	: data2 <= weights[1171];
				12'd1171	: data2 <= weights[1172];
				12'd1172	: data2 <= weights[1173];
				12'd1173	: data2 <= weights[1174];
				12'd1174	: data2 <= weights[1175];
				12'd1175	: data2 <= weights[1176];
				12'd1176	: data2 <= weights[1177];
				12'd1177	: data2 <= weights[1178];
				12'd1178	: data2 <= weights[1179];
				12'd1179	: data2 <= weights[1180];
				12'd1180	: data2 <= weights[1181];
				12'd1181	: data2 <= weights[1182];
				12'd1182	: data2 <= weights[1183];
				12'd1183	: data2 <= weights[1184];
				12'd1184	: data2 <= weights[1185];
				12'd1185	: data2 <= weights[1186];
				12'd1186	: data2 <= weights[1187];
				12'd1187	: data2 <= weights[1188];
				12'd1188	: data2 <= weights[1189];
				12'd1189	: data2 <= weights[1190];
				12'd1190	: data2 <= weights[1191];
				12'd1191	: data2 <= weights[1192];
				12'd1192	: data2 <= weights[1193];
				12'd1193	: data2 <= weights[1194];
				12'd1194	: data2 <= weights[1195];
				12'd1195	: data2 <= weights[1196];
				12'd1196	: data2 <= weights[1197];
				12'd1197	: data2 <= weights[1198];
				12'd1198	: data2 <= weights[1199];
				12'd1199	: data2 <= weights[1200];
				12'd1200	: data2 <= weights[1201];
				12'd1201	: data2 <= weights[1202];
				12'd1202	: data2 <= weights[1203];
				12'd1203	: data2 <= weights[1204];
				12'd1204	: data2 <= weights[1205];
				12'd1205	: data2 <= weights[1206];
				12'd1206	: data2 <= weights[1207];
				12'd1207	: data2 <= weights[1208];
				12'd1208	: data2 <= weights[1209];
				12'd1209	: data2 <= weights[1210];
				12'd1210	: data2 <= weights[1211];
				12'd1211	: data2 <= weights[1212];
				12'd1212	: data2 <= weights[1213];
				12'd1213	: data2 <= weights[1214];
				12'd1214	: data2 <= weights[1215];
				12'd1215	: data2 <= weights[1216];
				12'd1216	: data2 <= weights[1217];
				12'd1217	: data2 <= weights[1218];
				12'd1218	: data2 <= weights[1219];
				12'd1219	: data2 <= weights[1220];
				12'd1220	: data2 <= weights[1221];
				12'd1221	: data2 <= weights[1222];
				12'd1222	: data2 <= weights[1223];
				12'd1223	: data2 <= weights[1224];
				12'd1224	: data2 <= weights[1225];
				12'd1225	: data2 <= weights[1226];
				12'd1226	: data2 <= weights[1227];
				12'd1227	: data2 <= weights[1228];
				12'd1228	: data2 <= weights[1229];
				12'd1229	: data2 <= weights[1230];
				12'd1230	: data2 <= weights[1231];
				12'd1231	: data2 <= weights[1232];
				12'd1232	: data2 <= weights[1233];
				12'd1233	: data2 <= weights[1234];
				12'd1234	: data2 <= weights[1235];
				12'd1235	: data2 <= weights[1236];
				12'd1236	: data2 <= weights[1237];
				12'd1237	: data2 <= weights[1238];
				12'd1238	: data2 <= weights[1239];
				12'd1239	: data2 <= weights[1240];
				12'd1240	: data2 <= weights[1241];
				12'd1241	: data2 <= weights[1242];
				12'd1242	: data2 <= weights[1243];
				12'd1243	: data2 <= weights[1244];
				12'd1244	: data2 <= weights[1245];
				12'd1245	: data2 <= weights[1246];
				12'd1246	: data2 <= weights[1247];
				12'd1247	: data2 <= weights[1248];
				12'd1248	: data2 <= weights[1249];
				12'd1249	: data2 <= weights[1250];
				12'd1250	: data2 <= weights[1251];
				12'd1251	: data2 <= weights[1252];
				12'd1252	: data2 <= weights[1253];
				12'd1253	: data2 <= weights[1254];
				12'd1254	: data2 <= weights[1255];
				12'd1255	: data2 <= weights[1256];
				12'd1256	: data2 <= weights[1257];
				12'd1257	: data2 <= weights[1258];
				12'd1258	: data2 <= weights[1259];
				12'd1259	: data2 <= weights[1260];
				12'd1260	: data2 <= weights[1261];
				12'd1261	: data2 <= weights[1262];
				12'd1262	: data2 <= weights[1263];
				12'd1263	: data2 <= weights[1264];
				12'd1264	: data2 <= weights[1265];
				12'd1265	: data2 <= weights[1266];
				12'd1266	: data2 <= weights[1267];
				12'd1267	: data2 <= weights[1268];
				12'd1268	: data2 <= weights[1269];
				12'd1269	: data2 <= weights[1270];
				12'd1270	: data2 <= weights[1271];
				12'd1271	: data2 <= weights[1272];
				12'd1272	: data2 <= weights[1273];
				12'd1273	: data2 <= weights[1274];
				12'd1274	: data2 <= weights[1275];
				12'd1275	: data2 <= weights[1276];
				12'd1276	: data2 <= weights[1277];
				12'd1277	: data2 <= weights[1278];
				12'd1278	: data2 <= weights[1279];
				12'd1279	: data2 <= weights[1280];
				12'd1280	: data2 <= weights[1281];
				12'd1281	: data2 <= weights[1282];
				12'd1282	: data2 <= weights[1283];
				12'd1283	: data2 <= weights[1284];
				12'd1284	: data2 <= weights[1285];
				12'd1285	: data2 <= weights[1286];
				12'd1286	: data2 <= weights[1287];
				12'd1287	: data2 <= weights[1288];
				12'd1288	: data2 <= weights[1289];
				12'd1289	: data2 <= weights[1290];
				12'd1290	: data2 <= weights[1291];
				12'd1291	: data2 <= weights[1292];
				12'd1292	: data2 <= weights[1293];
				12'd1293	: data2 <= weights[1294];
				12'd1294	: data2 <= weights[1295];
				12'd1295	: data2 <= weights[1296];
				12'd1296	: data2 <= weights[1297];
				12'd1297	: data2 <= weights[1298];
				12'd1298	: data2 <= weights[1299];
				12'd1299	: data2 <= weights[1300];
				12'd1300	: data2 <= weights[1301];
				12'd1301	: data2 <= weights[1302];
				12'd1302	: data2 <= weights[1303];
				12'd1303	: data2 <= weights[1304];
				12'd1304	: data2 <= weights[1305];
				12'd1305	: data2 <= weights[1306];
				12'd1306	: data2 <= weights[1307];
				12'd1307	: data2 <= weights[1308];
				12'd1308	: data2 <= weights[1309];
				12'd1309	: data2 <= weights[1310];
				12'd1310	: data2 <= weights[1311];
				12'd1311	: data2 <= weights[1312];
				12'd1312	: data2 <= weights[1313];
				12'd1313	: data2 <= weights[1314];
				12'd1314	: data2 <= weights[1315];
				12'd1315	: data2 <= weights[1316];
				12'd1316	: data2 <= weights[1317];
				12'd1317	: data2 <= weights[1318];
				12'd1318	: data2 <= weights[1319];
				12'd1319	: data2 <= weights[1320];
				12'd1320	: data2 <= weights[1321];
				12'd1321	: data2 <= weights[1322];
				12'd1322	: data2 <= weights[1323];
				12'd1323	: data2 <= weights[1324];
				12'd1324	: data2 <= weights[1325];
				12'd1325	: data2 <= weights[1326];
				12'd1326	: data2 <= weights[1327];
				12'd1327	: data2 <= weights[1328];
				12'd1328	: data2 <= weights[1329];
				12'd1329	: data2 <= weights[1330];
				12'd1330	: data2 <= weights[1331];
				12'd1331	: data2 <= weights[1332];
				12'd1332	: data2 <= weights[1333];
				12'd1333	: data2 <= weights[1334];
				12'd1334	: data2 <= weights[1335];
				12'd1335	: data2 <= weights[1336];
				12'd1336	: data2 <= weights[1337];
				12'd1337	: data2 <= weights[1338];
				12'd1338	: data2 <= weights[1339];
				12'd1339	: data2 <= weights[1340];
				12'd1340	: data2 <= weights[1341];
				12'd1341	: data2 <= weights[1342];
				12'd1342	: data2 <= weights[1343];
				12'd1343	: data2 <= weights[1344];
				12'd1344	: data2 <= weights[1345];
				12'd1345	: data2 <= weights[1346];
				12'd1346	: data2 <= weights[1347];
				12'd1347	: data2 <= weights[1348];
				12'd1348	: data2 <= weights[1349];
				12'd1349	: data2 <= weights[1350];
				12'd1350	: data2 <= weights[1351];
				12'd1351	: data2 <= weights[1352];
				12'd1352	: data2 <= weights[1353];
				12'd1353	: data2 <= weights[1354];
				12'd1354	: data2 <= weights[1355];
				12'd1355	: data2 <= weights[1356];
				12'd1356	: data2 <= weights[1357];
				12'd1357	: data2 <= weights[1358];
				12'd1358	: data2 <= weights[1359];
				12'd1359	: data2 <= weights[1360];
				12'd1360	: data2 <= weights[1361];
				12'd1361	: data2 <= weights[1362];
				12'd1362	: data2 <= weights[1363];
				12'd1363	: data2 <= weights[1364];
				12'd1364	: data2 <= weights[1365];
				12'd1365	: data2 <= weights[1366];
				12'd1366	: data2 <= weights[1367];
				12'd1367	: data2 <= weights[1368];
				12'd1368	: data2 <= weights[1369];
				12'd1369	: data2 <= weights[1370];
				12'd1370	: data2 <= weights[1371];
				12'd1371	: data2 <= weights[1372];
				12'd1372	: data2 <= weights[1373];
				12'd1373	: data2 <= weights[1374];
				12'd1374	: data2 <= weights[1375];
				12'd1375	: data2 <= weights[1376];
				12'd1376	: data2 <= weights[1377];
				12'd1377	: data2 <= weights[1378];
				12'd1378	: data2 <= weights[1379];
				12'd1379	: data2 <= weights[1380];
				12'd1380	: data2 <= weights[1381];
				12'd1381	: data2 <= weights[1382];
				12'd1382	: data2 <= weights[1383];
				12'd1383	: data2 <= weights[1384];
				12'd1384	: data2 <= weights[1385];
				12'd1385	: data2 <= weights[1386];
				12'd1386	: data2 <= weights[1387];
				12'd1387	: data2 <= weights[1388];
				12'd1388	: data2 <= weights[1389];
				12'd1389	: data2 <= weights[1390];
				12'd1390	: data2 <= weights[1391];
				12'd1391	: data2 <= weights[1392];
				12'd1392	: data2 <= weights[1393];
				12'd1393	: data2 <= weights[1394];
				12'd1394	: data2 <= weights[1395];
				12'd1395	: data2 <= weights[1396];
				12'd1396	: data2 <= weights[1397];
				12'd1397	: data2 <= weights[1398];
				12'd1398	: data2 <= weights[1399];
				12'd1399	: data2 <= weights[1400];
				12'd1400	: data2 <= weights[1401];
				12'd1401	: data2 <= weights[1402];
				12'd1402	: data2 <= weights[1403];
				12'd1403	: data2 <= weights[1404];
				12'd1404	: data2 <= weights[1405];
				12'd1405	: data2 <= weights[1406];
				12'd1406	: data2 <= weights[1407];
				12'd1407	: data2 <= weights[1408];
				12'd1408	: data2 <= weights[1409];
				12'd1409	: data2 <= weights[1410];
				12'd1410	: data2 <= weights[1411];
				12'd1411	: data2 <= weights[1412];
				12'd1412	: data2 <= weights[1413];
				12'd1413	: data2 <= weights[1414];
				12'd1414	: data2 <= weights[1415];
				12'd1415	: data2 <= weights[1416];
				12'd1416	: data2 <= weights[1417];
				12'd1417	: data2 <= weights[1418];
				12'd1418	: data2 <= weights[1419];
				12'd1419	: data2 <= weights[1420];
				12'd1420	: data2 <= weights[1421];
				12'd1421	: data2 <= weights[1422];
				12'd1422	: data2 <= weights[1423];
				12'd1423	: data2 <= weights[1424];
				12'd1424	: data2 <= weights[1425];
				12'd1425	: data2 <= weights[1426];
				12'd1426	: data2 <= weights[1427];
				12'd1427	: data2 <= weights[1428];
				12'd1428	: data2 <= weights[1429];
				12'd1429	: data2 <= weights[1430];
				12'd1430	: data2 <= weights[1431];
				12'd1431	: data2 <= weights[1432];
				12'd1432	: data2 <= weights[1433];
				12'd1433	: data2 <= weights[1434];
				12'd1434	: data2 <= weights[1435];
				12'd1435	: data2 <= weights[1436];
				12'd1436	: data2 <= weights[1437];
				12'd1437	: data2 <= weights[1438];
				12'd1438	: data2 <= weights[1439];
				12'd1439	: data2 <= weights[1440];
				12'd1440	: data2 <= weights[1441];
				12'd1441	: data2 <= weights[1442];
				12'd1442	: data2 <= weights[1443];
				12'd1443	: data2 <= weights[1444];
				12'd1444	: data2 <= weights[1445];
				12'd1445	: data2 <= weights[1446];
				12'd1446	: data2 <= weights[1447];
				12'd1447	: data2 <= weights[1448];
				12'd1448	: data2 <= weights[1449];
				12'd1449	: data2 <= weights[1450];
				12'd1450	: data2 <= weights[1451];
				12'd1451	: data2 <= weights[1452];
				12'd1452	: data2 <= weights[1453];
				12'd1453	: data2 <= weights[1454];
				12'd1454	: data2 <= weights[1455];
				12'd1455	: data2 <= weights[1456];
				12'd1456	: data2 <= weights[1457];
				12'd1457	: data2 <= weights[1458];
				12'd1458	: data2 <= weights[1459];
				12'd1459	: data2 <= weights[1460];
				12'd1460	: data2 <= weights[1461];
				12'd1461	: data2 <= weights[1462];
				12'd1462	: data2 <= weights[1463];
				12'd1463	: data2 <= weights[1464];
				12'd1464	: data2 <= weights[1465];
				12'd1465	: data2 <= weights[1466];
				12'd1466	: data2 <= weights[1467];
				12'd1467	: data2 <= weights[1468];
				12'd1468	: data2 <= weights[1469];
				12'd1469	: data2 <= weights[1470];
				12'd1470	: data2 <= weights[1471];
				12'd1471	: data2 <= weights[1472];
				12'd1472	: data2 <= weights[1473];
				12'd1473	: data2 <= weights[1474];
				12'd1474	: data2 <= weights[1475];
				12'd1475	: data2 <= weights[1476];
				12'd1476	: data2 <= weights[1477];
				12'd1477	: data2 <= weights[1478];
				12'd1478	: data2 <= weights[1479];
				12'd1479	: data2 <= weights[1480];
				12'd1480	: data2 <= weights[1481];
				12'd1481	: data2 <= weights[1482];
				12'd1482	: data2 <= weights[1483];
				12'd1483	: data2 <= weights[1484];
				12'd1484	: data2 <= weights[1485];
				12'd1485	: data2 <= weights[1486];
				12'd1486	: data2 <= weights[1487];
				12'd1487	: data2 <= weights[1488];
				12'd1488	: data2 <= weights[1489];
				12'd1489	: data2 <= weights[1490];
				12'd1490	: data2 <= weights[1491];
				12'd1491	: data2 <= weights[1492];
				12'd1492	: data2 <= weights[1493];
				12'd1493	: data2 <= weights[1494];
				12'd1494	: data2 <= weights[1495];
				12'd1495	: data2 <= weights[1496];
				12'd1496	: data2 <= weights[1497];
				12'd1497	: data2 <= weights[1498];
				12'd1498	: data2 <= weights[1499];
				12'd1499	: data2 <= weights[1500];
				12'd1500	: data2 <= weights[1501];
				12'd1501	: data2 <= weights[1502];
				12'd1502	: data2 <= weights[1503];
				12'd1503	: data2 <= weights[1504];
				12'd1504	: data2 <= weights[1505];
				12'd1505	: data2 <= weights[1506];
				12'd1506	: data2 <= weights[1507];
				12'd1507	: data2 <= weights[1508];
				12'd1508	: data2 <= weights[1509];
				12'd1509	: data2 <= weights[1510];
				12'd1510	: data2 <= weights[1511];
				12'd1511	: data2 <= weights[1512];
				12'd1512	: data2 <= weights[1513];
				12'd1513	: data2 <= weights[1514];
				12'd1514	: data2 <= weights[1515];
				12'd1515	: data2 <= weights[1516];
				12'd1516	: data2 <= weights[1517];
				12'd1517	: data2 <= weights[1518];
				12'd1518	: data2 <= weights[1519];
				12'd1519	: data2 <= weights[1520];
				12'd1520	: data2 <= weights[1521];
				12'd1521	: data2 <= weights[1522];
				12'd1522	: data2 <= weights[1523];
				12'd1523	: data2 <= weights[1524];
				12'd1524	: data2 <= weights[1525];
				12'd1525	: data2 <= weights[1526];
				12'd1526	: data2 <= weights[1527];
				12'd1527	: data2 <= weights[1528];
				12'd1528	: data2 <= weights[1529];
				12'd1529	: data2 <= weights[1530];
				12'd1530	: data2 <= weights[1531];
				12'd1531	: data2 <= weights[1532];
				12'd1532	: data2 <= weights[1533];
				12'd1533	: data2 <= weights[1534];
				12'd1534	: data2 <= weights[1535];
				12'd1535	: data2 <= weights[1536];
				12'd1536	: data2 <= weights[1537];
				12'd1537	: data2 <= weights[1538];
				12'd1538	: data2 <= weights[1539];
				12'd1539	: data2 <= weights[1540];
				12'd1540	: data2 <= weights[1541];
				12'd1541	: data2 <= weights[1542];
				12'd1542	: data2 <= weights[1543];
				12'd1543	: data2 <= weights[1544];
				12'd1544	: data2 <= weights[1545];
				12'd1545	: data2 <= weights[1546];
				12'd1546	: data2 <= weights[1547];
				12'd1547	: data2 <= weights[1548];
				12'd1548	: data2 <= weights[1549];
				12'd1549	: data2 <= weights[1550];
				12'd1550	: data2 <= weights[1551];
				12'd1551	: data2 <= weights[1552];
				12'd1552	: data2 <= weights[1553];
				12'd1553	: data2 <= weights[1554];
				12'd1554	: data2 <= weights[1555];
				12'd1555	: data2 <= weights[1556];
				12'd1556	: data2 <= weights[1557];
				12'd1557	: data2 <= weights[1558];
				12'd1558	: data2 <= weights[1559];
				12'd1559	: data2 <= weights[1560];
				12'd1560	: data2 <= weights[1561];
				12'd1561	: data2 <= weights[1562];
				12'd1562	: data2 <= weights[1563];
				12'd1563	: data2 <= weights[1564];
				12'd1564	: data2 <= weights[1565];
				12'd1565	: data2 <= weights[1566];
				12'd1566	: data2 <= weights[1567];
				12'd1567	: data2 <= weights[1568];
				12'd1568	: data2 <= weights[1569];
				12'd1569	: data2 <= weights[1570];
				12'd1570	: data2 <= weights[1571];
				12'd1571	: data2 <= weights[1572];
				12'd1572	: data2 <= weights[1573];
				12'd1573	: data2 <= weights[1574];
				12'd1574	: data2 <= weights[1575];
				12'd1575	: data2 <= weights[1576];
				12'd1576	: data2 <= weights[1577];
				12'd1577	: data2 <= weights[1578];
				12'd1578	: data2 <= weights[1579];
				12'd1579	: data2 <= weights[1580];
				12'd1580	: data2 <= weights[1581];
				12'd1581	: data2 <= weights[1582];
				12'd1582	: data2 <= weights[1583];
				12'd1583	: data2 <= weights[1584];
				12'd1584	: data2 <= weights[1585];
				12'd1585	: data2 <= weights[1586];
				12'd1586	: data2 <= weights[1587];
				12'd1587	: data2 <= weights[1588];
				12'd1588	: data2 <= weights[1589];
				12'd1589	: data2 <= weights[1590];
				12'd1590	: data2 <= weights[1591];
				12'd1591	: data2 <= weights[1592];
				12'd1592	: data2 <= weights[1593];
				12'd1593	: data2 <= weights[1594];
				12'd1594	: data2 <= weights[1595];
				12'd1595	: data2 <= weights[1596];
				12'd1596	: data2 <= weights[1597];
				12'd1597	: data2 <= weights[1598];
				12'd1598	: data2 <= weights[1599];
				12'd1599	: data2 <= weights[1600];
				12'd1600	: data2 <= weights[1601];
				12'd1601	: data2 <= weights[1602];
				12'd1602	: data2 <= weights[1603];
				12'd1603	: data2 <= weights[1604];
				12'd1604	: data2 <= weights[1605];
				12'd1605	: data2 <= weights[1606];
				12'd1606	: data2 <= weights[1607];
				12'd1607	: data2 <= weights[1608];
				12'd1608	: data2 <= weights[1609];
				12'd1609	: data2 <= weights[1610];
				12'd1610	: data2 <= weights[1611];
				12'd1611	: data2 <= weights[1612];
				12'd1612	: data2 <= weights[1613];
				12'd1613	: data2 <= weights[1614];
				12'd1614	: data2 <= weights[1615];
				12'd1615	: data2 <= weights[1616];
				12'd1616	: data2 <= weights[1617];
				12'd1617	: data2 <= weights[1618];
				12'd1618	: data2 <= weights[1619];
				12'd1619	: data2 <= weights[1620];
				12'd1620	: data2 <= weights[1621];
				12'd1621	: data2 <= weights[1622];
				12'd1622	: data2 <= weights[1623];
				12'd1623	: data2 <= weights[1624];
				12'd1624	: data2 <= weights[1625];
				12'd1625	: data2 <= weights[1626];
				12'd1626	: data2 <= weights[1627];
				12'd1627	: data2 <= weights[1628];
				12'd1628	: data2 <= weights[1629];
				12'd1629	: data2 <= weights[1630];
				12'd1630	: data2 <= weights[1631];
				12'd1631	: data2 <= weights[1632];
				12'd1632	: data2 <= weights[1633];
				12'd1633	: data2 <= weights[1634];
				12'd1634	: data2 <= weights[1635];
				12'd1635	: data2 <= weights[1636];
				12'd1636	: data2 <= weights[1637];
				12'd1637	: data2 <= weights[1638];
				12'd1638	: data2 <= weights[1639];
				12'd1639	: data2 <= weights[1640];
				12'd1640	: data2 <= weights[1641];
				12'd1641	: data2 <= weights[1642];
				12'd1642	: data2 <= weights[1643];
				12'd1643	: data2 <= weights[1644];
				12'd1644	: data2 <= weights[1645];
				12'd1645	: data2 <= weights[1646];
				12'd1646	: data2 <= weights[1647];
				12'd1647	: data2 <= weights[1648];
				12'd1648	: data2 <= weights[1649];
				12'd1649	: data2 <= weights[1650];
				12'd1650	: data2 <= weights[1651];
				12'd1651	: data2 <= weights[1652];
				12'd1652	: data2 <= weights[1653];
				12'd1653	: data2 <= weights[1654];
				12'd1654	: data2 <= weights[1655];
				12'd1655	: data2 <= weights[1656];
				12'd1656	: data2 <= weights[1657];
				12'd1657	: data2 <= weights[1658];
				12'd1658	: data2 <= weights[1659];
				12'd1659	: data2 <= weights[1660];
				12'd1660	: data2 <= weights[1661];
				12'd1661	: data2 <= weights[1662];
				12'd1662	: data2 <= weights[1663];
				12'd1663	: data2 <= weights[1664];
				12'd1664	: data2 <= weights[1665];
				12'd1665	: data2 <= weights[1666];
				12'd1666	: data2 <= weights[1667];
				12'd1667	: data2 <= weights[1668];
				12'd1668	: data2 <= weights[1669];
				12'd1669	: data2 <= weights[1670];
				12'd1670	: data2 <= weights[1671];
				12'd1671	: data2 <= weights[1672];
				12'd1672	: data2 <= weights[1673];
				12'd1673	: data2 <= weights[1674];
				12'd1674	: data2 <= weights[1675];
				12'd1675	: data2 <= weights[1676];
				12'd1676	: data2 <= weights[1677];
				12'd1677	: data2 <= weights[1678];
				12'd1678	: data2 <= weights[1679];
				12'd1679	: data2 <= weights[1680];
				12'd1680	: data2 <= weights[1681];
				12'd1681	: data2 <= weights[1682];
				12'd1682	: data2 <= weights[1683];
				12'd1683	: data2 <= weights[1684];
				12'd1684	: data2 <= weights[1685];
				12'd1685	: data2 <= weights[1686];
				12'd1686	: data2 <= weights[1687];
				12'd1687	: data2 <= weights[1688];
				12'd1688	: data2 <= weights[1689];
				12'd1689	: data2 <= weights[1690];
				12'd1690	: data2 <= weights[1691];
				12'd1691	: data2 <= weights[1692];
				12'd1692	: data2 <= weights[1693];
				12'd1693	: data2 <= weights[1694];
				12'd1694	: data2 <= weights[1695];
				12'd1695	: data2 <= weights[1696];
				12'd1696	: data2 <= weights[1697];
				12'd1697	: data2 <= weights[1698];
				12'd1698	: data2 <= weights[1699];
				12'd1699	: data2 <= weights[1700];
				12'd1700	: data2 <= weights[1701];
				12'd1701	: data2 <= weights[1702];
				12'd1702	: data2 <= weights[1703];
				12'd1703	: data2 <= weights[1704];
				12'd1704	: data2 <= weights[1705];
				12'd1705	: data2 <= weights[1706];
				12'd1706	: data2 <= weights[1707];
				12'd1707	: data2 <= weights[1708];
				12'd1708	: data2 <= weights[1709];
				12'd1709	: data2 <= weights[1710];
				12'd1710	: data2 <= weights[1711];
				12'd1711	: data2 <= weights[1712];
				12'd1712	: data2 <= weights[1713];
				12'd1713	: data2 <= weights[1714];
				12'd1714	: data2 <= weights[1715];
				12'd1715	: data2 <= weights[1716];
				12'd1716	: data2 <= weights[1717];
				12'd1717	: data2 <= weights[1718];
				12'd1718	: data2 <= weights[1719];
				12'd1719	: data2 <= weights[1720];
				12'd1720	: data2 <= weights[1721];
				12'd1721	: data2 <= weights[1722];
				12'd1722	: data2 <= weights[1723];
				12'd1723	: data2 <= weights[1724];
				12'd1724	: data2 <= weights[1725];
				12'd1725	: data2 <= weights[1726];
				12'd1726	: data2 <= weights[1727];
				12'd1727	: data2 <= weights[1728];
				12'd1728	: data2 <= weights[1729];
				12'd1729	: data2 <= weights[1730];
				12'd1730	: data2 <= weights[1731];
				12'd1731	: data2 <= weights[1732];
				12'd1732	: data2 <= weights[1733];
				12'd1733	: data2 <= weights[1734];
				12'd1734	: data2 <= weights[1735];
				12'd1735	: data2 <= weights[1736];
				12'd1736	: data2 <= weights[1737];
				12'd1737	: data2 <= weights[1738];
				12'd1738	: data2 <= weights[1739];
				12'd1739	: data2 <= weights[1740];
				12'd1740	: data2 <= weights[1741];
				12'd1741	: data2 <= weights[1742];
				12'd1742	: data2 <= weights[1743];
				12'd1743	: data2 <= weights[1744];
				12'd1744	: data2 <= weights[1745];
				12'd1745	: data2 <= weights[1746];
				12'd1746	: data2 <= weights[1747];
				12'd1747	: data2 <= weights[1748];
				12'd1748	: data2 <= weights[1749];
				12'd1749	: data2 <= weights[1750];
				12'd1750	: data2 <= weights[1751];
				12'd1751	: data2 <= weights[1752];
				12'd1752	: data2 <= weights[1753];
				12'd1753	: data2 <= weights[1754];
				12'd1754	: data2 <= weights[1755];
				12'd1755	: data2 <= weights[1756];
				12'd1756	: data2 <= weights[1757];
				12'd1757	: data2 <= weights[1758];
				12'd1758	: data2 <= weights[1759];
				12'd1759	: data2 <= weights[1760];
				12'd1760	: data2 <= weights[1761];
				12'd1761	: data2 <= weights[1762];
				12'd1762	: data2 <= weights[1763];
				12'd1763	: data2 <= weights[1764];
				12'd1764	: data2 <= weights[1765];
				12'd1765	: data2 <= weights[1766];
				12'd1766	: data2 <= weights[1767];
				12'd1767	: data2 <= weights[1768];
				12'd1768	: data2 <= weights[1769];
				12'd1769	: data2 <= weights[1770];
				12'd1770	: data2 <= weights[1771];
				12'd1771	: data2 <= weights[1772];
				12'd1772	: data2 <= weights[1773];
				12'd1773	: data2 <= weights[1774];
				12'd1774	: data2 <= weights[1775];
				12'd1775	: data2 <= weights[1776];
				12'd1776	: data2 <= weights[1777];
				12'd1777	: data2 <= weights[1778];
				12'd1778	: data2 <= weights[1779];
				12'd1779	: data2 <= weights[1780];
				12'd1780	: data2 <= weights[1781];
				12'd1781	: data2 <= weights[1782];
				12'd1782	: data2 <= weights[1783];
				12'd1783	: data2 <= weights[1784];
				12'd1784	: data2 <= weights[1785];
				12'd1785	: data2 <= weights[1786];
				12'd1786	: data2 <= weights[1787];
				12'd1787	: data2 <= weights[1788];
				12'd1788	: data2 <= weights[1789];
				12'd1789	: data2 <= weights[1790];
				12'd1790	: data2 <= weights[1791];
				12'd1791	: data2 <= weights[1792];
				12'd1792	: data2 <= weights[1793];
				12'd1793	: data2 <= weights[1794];
				12'd1794	: data2 <= weights[1795];
				12'd1795	: data2 <= weights[1796];
				12'd1796	: data2 <= weights[1797];
				12'd1797	: data2 <= weights[1798];
				12'd1798	: data2 <= weights[1799];
				12'd1799	: data2 <= weights[1800];
				12'd1800	: data2 <= weights[1801];
				12'd1801	: data2 <= weights[1802];
				12'd1802	: data2 <= weights[1803];
				12'd1803	: data2 <= weights[1804];
				12'd1804	: data2 <= weights[1805];
				12'd1805	: data2 <= weights[1806];
				12'd1806	: data2 <= weights[1807];
				12'd1807	: data2 <= weights[1808];
				12'd1808	: data2 <= weights[1809];
				12'd1809	: data2 <= weights[1810];
				12'd1810	: data2 <= weights[1811];
				12'd1811	: data2 <= weights[1812];
				12'd1812	: data2 <= weights[1813];
				12'd1813	: data2 <= weights[1814];
				12'd1814	: data2 <= weights[1815];
				12'd1815	: data2 <= weights[1816];
				12'd1816	: data2 <= weights[1817];
				12'd1817	: data2 <= weights[1818];
				12'd1818	: data2 <= weights[1819];
				12'd1819	: data2 <= weights[1820];
				12'd1820	: data2 <= weights[1821];
				12'd1821	: data2 <= weights[1822];
				12'd1822	: data2 <= weights[1823];
				12'd1823	: data2 <= weights[1824];
				12'd1824	: data2 <= weights[1825];
				12'd1825	: data2 <= weights[1826];
				12'd1826	: data2 <= weights[1827];
				12'd1827	: data2 <= weights[1828];
				12'd1828	: data2 <= weights[1829];
				12'd1829	: data2 <= weights[1830];
				12'd1830	: data2 <= weights[1831];
				12'd1831	: data2 <= weights[1832];
				12'd1832	: data2 <= weights[1833];
				12'd1833	: data2 <= weights[1834];
				12'd1834	: data2 <= weights[1835];
				12'd1835	: data2 <= weights[1836];
				12'd1836	: data2 <= weights[1837];
				12'd1837	: data2 <= weights[1838];
				12'd1838	: data2 <= weights[1839];
				12'd1839	: data2 <= weights[1840];
				12'd1840	: data2 <= weights[1841];
				12'd1841	: data2 <= weights[1842];
				12'd1842	: data2 <= weights[1843];
				12'd1843	: data2 <= weights[1844];
				12'd1844	: data2 <= weights[1845];
				12'd1845	: data2 <= weights[1846];
				12'd1846	: data2 <= weights[1847];
				12'd1847	: data2 <= weights[1848];
				12'd1848	: data2 <= weights[1849];
				12'd1849	: data2 <= weights[1850];
				12'd1850	: data2 <= weights[1851];
				12'd1851	: data2 <= weights[1852];
				12'd1852	: data2 <= weights[1853];
				12'd1853	: data2 <= weights[1854];
				12'd1854	: data2 <= weights[1855];
				12'd1855	: data2 <= weights[1856];
				12'd1856	: data2 <= weights[1857];
				12'd1857	: data2 <= weights[1858];
				12'd1858	: data2 <= weights[1859];
				12'd1859	: data2 <= weights[1860];
				12'd1860	: data2 <= weights[1861];
				12'd1861	: data2 <= weights[1862];
				12'd1862	: data2 <= weights[1863];
				12'd1863	: data2 <= weights[1864];
				12'd1864	: data2 <= weights[1865];
				12'd1865	: data2 <= weights[1866];
				12'd1866	: data2 <= weights[1867];
				12'd1867	: data2 <= weights[1868];
				12'd1868	: data2 <= weights[1869];
				12'd1869	: data2 <= weights[1870];
				12'd1870	: data2 <= weights[1871];
				12'd1871	: data2 <= weights[1872];
				12'd1872	: data2 <= weights[1873];
				12'd1873	: data2 <= weights[1874];
				12'd1874	: data2 <= weights[1875];
				12'd1875	: data2 <= weights[1876];
				12'd1876	: data2 <= weights[1877];
				12'd1877	: data2 <= weights[1878];
				12'd1878	: data2 <= weights[1879];
				12'd1879	: data2 <= weights[1880];
				12'd1880	: data2 <= weights[1881];
				12'd1881	: data2 <= weights[1882];
				12'd1882	: data2 <= weights[1883];
				12'd1883	: data2 <= weights[1884];
				12'd1884	: data2 <= weights[1885];
				12'd1885	: data2 <= weights[1886];
				12'd1886	: data2 <= weights[1887];
				12'd1887	: data2 <= weights[1888];
				12'd1888	: data2 <= weights[1889];
				12'd1889	: data2 <= weights[1890];
				12'd1890	: data2 <= weights[1891];
				12'd1891	: data2 <= weights[1892];
				12'd1892	: data2 <= weights[1893];
				12'd1893	: data2 <= weights[1894];
				12'd1894	: data2 <= weights[1895];
				12'd1895	: data2 <= weights[1896];
				12'd1896	: data2 <= weights[1897];
				12'd1897	: data2 <= weights[1898];
				12'd1898	: data2 <= weights[1899];
				12'd1899	: data2 <= weights[1900];
				12'd1900	: data2 <= weights[1901];
				12'd1901	: data2 <= weights[1902];
				12'd1902	: data2 <= weights[1903];
				12'd1903	: data2 <= weights[1904];
				12'd1904	: data2 <= weights[1905];
				12'd1905	: data2 <= weights[1906];
				12'd1906	: data2 <= weights[1907];
				12'd1907	: data2 <= weights[1908];
				12'd1908	: data2 <= weights[1909];
				12'd1909	: data2 <= weights[1910];
				12'd1910	: data2 <= weights[1911];
				12'd1911	: data2 <= weights[1912];
				12'd1912	: data2 <= weights[1913];
				12'd1913	: data2 <= weights[1914];
				12'd1914	: data2 <= weights[1915];
				12'd1915	: data2 <= weights[1916];
				12'd1916	: data2 <= weights[1917];
				12'd1917	: data2 <= weights[1918];
				12'd1918	: data2 <= weights[1919];
				12'd1919	: data2 <= weights[1920];
				12'd1920	: data2 <= weights[1921];
				12'd1921	: data2 <= weights[1922];
				12'd1922	: data2 <= weights[1923];
				12'd1923	: data2 <= weights[1924];
				12'd1924	: data2 <= weights[1925];
				12'd1925	: data2 <= weights[1926];
				12'd1926	: data2 <= weights[1927];
				12'd1927	: data2 <= weights[1928];
				12'd1928	: data2 <= weights[1929];
				12'd1929	: data2 <= weights[1930];
				12'd1930	: data2 <= weights[1931];
				12'd1931	: data2 <= weights[1932];
				12'd1932	: data2 <= weights[1933];
				12'd1933	: data2 <= weights[1934];
				12'd1934	: data2 <= weights[1935];
				12'd1935	: data2 <= weights[1936];
				12'd1936	: data2 <= weights[1937];
				12'd1937	: data2 <= weights[1938];
				12'd1938	: data2 <= weights[1939];
				12'd1939	: data2 <= weights[1940];
				12'd1940	: data2 <= weights[1941];
				12'd1941	: data2 <= weights[1942];
				12'd1942	: data2 <= weights[1943];
				12'd1943	: data2 <= weights[1944];
				12'd1944	: data2 <= weights[1945];
				12'd1945	: data2 <= weights[1946];
				12'd1946	: data2 <= weights[1947];
				12'd1947	: data2 <= weights[1948];
				12'd1948	: data2 <= weights[1949];
				12'd1949	: data2 <= weights[1950];
				12'd1950	: data2 <= weights[1951];
				12'd1951	: data2 <= weights[1952];
				12'd1952	: data2 <= weights[1953];
				12'd1953	: data2 <= weights[1954];
				12'd1954	: data2 <= weights[1955];
				12'd1955	: data2 <= weights[1956];
				12'd1956	: data2 <= weights[1957];
				12'd1957	: data2 <= weights[1958];
				12'd1958	: data2 <= weights[1959];
				12'd1959	: data2 <= weights[1960];
				12'd1960	: data2 <= weights[1961];
				12'd1961	: data2 <= weights[1962];
				12'd1962	: data2 <= weights[1963];
				12'd1963	: data2 <= weights[1964];
				12'd1964	: data2 <= weights[1965];
				12'd1965	: data2 <= weights[1966];
				12'd1966	: data2 <= weights[1967];
				12'd1967	: data2 <= weights[1968];
				12'd1968	: data2 <= weights[1969];
				12'd1969	: data2 <= weights[1970];
				12'd1970	: data2 <= weights[1971];
				12'd1971	: data2 <= weights[1972];
				12'd1972	: data2 <= weights[1973];
				12'd1973	: data2 <= weights[1974];
				12'd1974	: data2 <= weights[1975];
				12'd1975	: data2 <= weights[1976];
				12'd1976	: data2 <= weights[1977];
				12'd1977	: data2 <= weights[1978];
				12'd1978	: data2 <= weights[1979];
				12'd1979	: data2 <= weights[1980];
				12'd1980	: data2 <= weights[1981];
				12'd1981	: data2 <= weights[1982];
				12'd1982	: data2 <= weights[1983];
				12'd1983	: data2 <= weights[1984];
				12'd1984	: data2 <= weights[1985];
				12'd1985	: data2 <= weights[1986];
				12'd1986	: data2 <= weights[1987];
				12'd1987	: data2 <= weights[1988];
				12'd1988	: data2 <= weights[1989];
				12'd1989	: data2 <= weights[1990];
				12'd1990	: data2 <= weights[1991];
				12'd1991	: data2 <= weights[1992];
				12'd1992	: data2 <= weights[1993];
				12'd1993	: data2 <= weights[1994];
				12'd1994	: data2 <= weights[1995];
				12'd1995	: data2 <= weights[1996];
				12'd1996	: data2 <= weights[1997];
				12'd1997	: data2 <= weights[1998];
				12'd1998	: data2 <= weights[1999];
				12'd1999	: data2 <= weights[2000];
				12'd2000	: data2 <= weights[2001];
				12'd2001	: data2 <= weights[2002];
				12'd2002	: data2 <= weights[2003];
				12'd2003	: data2 <= weights[2004];
				12'd2004	: data2 <= weights[2005];
				12'd2005	: data2 <= weights[2006];
				12'd2006	: data2 <= weights[2007];
				12'd2007	: data2 <= weights[2008];
				12'd2008	: data2 <= weights[2009];
				12'd2009	: data2 <= weights[2010];
				12'd2010	: data2 <= weights[2011];
				12'd2011	: data2 <= weights[2012];
				12'd2012	: data2 <= weights[2013];
				12'd2013	: data2 <= weights[2014];
				12'd2014	: data2 <= weights[2015];
				12'd2015	: data2 <= weights[2016];
				12'd2016	: data2 <= weights[2017];
				12'd2017	: data2 <= weights[2018];
				12'd2018	: data2 <= weights[2019];
				12'd2019	: data2 <= weights[2020];
				12'd2020	: data2 <= weights[2021];
				12'd2021	: data2 <= weights[2022];
				12'd2022	: data2 <= weights[2023];
				12'd2023	: data2 <= weights[2024];
				12'd2024	: data2 <= weights[2025];
				12'd2025	: data2 <= weights[2026];
				12'd2026	: data2 <= weights[2027];
				12'd2027	: data2 <= weights[2028];
				12'd2028	: data2 <= weights[2029];
				12'd2029	: data2 <= weights[2030];
				12'd2030	: data2 <= weights[2031];
				12'd2031	: data2 <= weights[2032];
				12'd2032	: data2 <= weights[2033];
				12'd2033	: data2 <= weights[2034];
				12'd2034	: data2 <= weights[2035];
				12'd2035	: data2 <= weights[2036];
				12'd2036	: data2 <= weights[2037];
				12'd2037	: data2 <= weights[2038];
				12'd2038	: data2 <= weights[2039];
				12'd2039	: data2 <= weights[2040];
				12'd2040	: data2 <= weights[2041];
				12'd2041	: data2 <= weights[2042];
				12'd2042	: data2 <= weights[2043];
				12'd2043	: data2 <= weights[2044];
				12'd2044	: data2 <= weights[2045];
				12'd2045	: data2 <= weights[2046];
				12'd2046	: data2 <= weights[2047];
				12'd2047	: data2 <= weights[2048];
				12'd2048	: data2 <= weights[2049];
				12'd2049	: data2 <= weights[2050];
				12'd2050	: data2 <= weights[2051];
				12'd2051	: data2 <= weights[2052];
				12'd2052	: data2 <= weights[2053];
				12'd2053	: data2 <= weights[2054];
				12'd2054	: data2 <= weights[2055];
				12'd2055	: data2 <= weights[2056];
				12'd2056	: data2 <= weights[2057];
				12'd2057	: data2 <= weights[2058];
				12'd2058	: data2 <= weights[2059];
				12'd2059	: data2 <= weights[2060];
				12'd2060	: data2 <= weights[2061];
				12'd2061	: data2 <= weights[2062];
				12'd2062	: data2 <= weights[2063];
				12'd2063	: data2 <= weights[2064];
				12'd2064	: data2 <= weights[2065];
				12'd2065	: data2 <= weights[2066];
				12'd2066	: data2 <= weights[2067];
				12'd2067	: data2 <= weights[2068];
				12'd2068	: data2 <= weights[2069];
				12'd2069	: data2 <= weights[2070];
				12'd2070	: data2 <= weights[2071];
				12'd2071	: data2 <= weights[2072];
				12'd2072	: data2 <= weights[2073];
				12'd2073	: data2 <= weights[2074];
				12'd2074	: data2 <= weights[2075];
				12'd2075	: data2 <= weights[2076];
				12'd2076	: data2 <= weights[2077];
				12'd2077	: data2 <= weights[2078];
				12'd2078	: data2 <= weights[2079];
				12'd2079	: data2 <= weights[2080];
				12'd2080	: data2 <= weights[2081];
				12'd2081	: data2 <= weights[2082];
				12'd2082	: data2 <= weights[2083];
				12'd2083	: data2 <= weights[2084];
				12'd2084	: data2 <= weights[2085];
				12'd2085	: data2 <= weights[2086];
				12'd2086	: data2 <= weights[2087];
				12'd2087	: data2 <= weights[2088];
				12'd2088	: data2 <= weights[2089];
				12'd2089	: data2 <= weights[2090];
				12'd2090	: data2 <= weights[2091];
				12'd2091	: data2 <= weights[2092];
				12'd2092	: data2 <= weights[2093];
				12'd2093	: data2 <= weights[2094];
				12'd2094	: data2 <= weights[2095];
				12'd2095	: data2 <= weights[2096];
				12'd2096	: data2 <= weights[2097];
				12'd2097	: data2 <= weights[2098];
				12'd2098	: data2 <= weights[2099];
				12'd2099	: data2 <= weights[2100];
				12'd2100	: data2 <= weights[2101];
				12'd2101	: data2 <= weights[2102];
				12'd2102	: data2 <= weights[2103];
				12'd2103	: data2 <= weights[2104];
				12'd2104	: data2 <= weights[2105];
				12'd2105	: data2 <= weights[2106];
				12'd2106	: data2 <= weights[2107];
				12'd2107	: data2 <= weights[2108];
				12'd2108	: data2 <= weights[2109];
				12'd2109	: data2 <= weights[2110];
				12'd2110	: data2 <= weights[2111];
				12'd2111	: data2 <= weights[2112];
				12'd2112	: data2 <= weights[2113];
				12'd2113	: data2 <= weights[2114];
				12'd2114	: data2 <= weights[2115];
				12'd2115	: data2 <= weights[2116];
				12'd2116	: data2 <= weights[2117];
				12'd2117	: data2 <= weights[2118];
				12'd2118	: data2 <= weights[2119];
				12'd2119	: data2 <= weights[2120];
				12'd2120	: data2 <= weights[2121];
				12'd2121	: data2 <= weights[2122];
				12'd2122	: data2 <= weights[2123];
				12'd2123	: data2 <= weights[2124];
				12'd2124	: data2 <= weights[2125];
				12'd2125	: data2 <= weights[2126];
				12'd2126	: data2 <= weights[2127];
				12'd2127	: data2 <= weights[2128];
				12'd2128	: data2 <= weights[2129];
				12'd2129	: data2 <= weights[2130];
				12'd2130	: data2 <= weights[2131];
				12'd2131	: data2 <= weights[2132];
				12'd2132	: data2 <= weights[2133];
				12'd2133	: data2 <= weights[2134];
				12'd2134	: data2 <= weights[2135];
				12'd2135	: data2 <= weights[2136];
				12'd2136	: data2 <= weights[2137];
				12'd2137	: data2 <= weights[2138];
				12'd2138	: data2 <= weights[2139];
				12'd2139	: data2 <= weights[2140];
				12'd2140	: data2 <= weights[2141];
				12'd2141	: data2 <= weights[2142];
				12'd2142	: data2 <= weights[2143];
				12'd2143	: data2 <= weights[2144];
				12'd2144	: data2 <= weights[2145];
				12'd2145	: data2 <= weights[2146];
				12'd2146	: data2 <= weights[2147];
				12'd2147	: data2 <= weights[2148];
				12'd2148	: data2 <= weights[2149];
				12'd2149	: data2 <= weights[2150];
				12'd2150	: data2 <= weights[2151];
				12'd2151	: data2 <= weights[2152];
				12'd2152	: data2 <= weights[2153];
				12'd2153	: data2 <= weights[2154];
				12'd2154	: data2 <= weights[2155];
				12'd2155	: data2 <= weights[2156];
				12'd2156	: data2 <= weights[2157];
				12'd2157	: data2 <= weights[2158];
				12'd2158	: data2 <= weights[2159];
				12'd2159	: data2 <= weights[2160];
				12'd2160	: data2 <= weights[2161];
				12'd2161	: data2 <= weights[2162];
				12'd2162	: data2 <= weights[2163];
				12'd2163	: data2 <= weights[2164];
				12'd2164	: data2 <= weights[2165];
				12'd2165	: data2 <= weights[2166];
				12'd2166	: data2 <= weights[2167];
				12'd2167	: data2 <= weights[2168];
				12'd2168	: data2 <= weights[2169];
				12'd2169	: data2 <= weights[2170];
				12'd2170	: data2 <= weights[2171];
				12'd2171	: data2 <= weights[2172];
				12'd2172	: data2 <= weights[2173];
				12'd2173	: data2 <= weights[2174];
				12'd2174	: data2 <= weights[2175];
				12'd2175	: data2 <= weights[2176];
				12'd2176	: data2 <= weights[2177];
				12'd2177	: data2 <= weights[2178];
				12'd2178	: data2 <= weights[2179];
				12'd2179	: data2 <= weights[2180];
				12'd2180	: data2 <= weights[2181];
				12'd2181	: data2 <= weights[2182];
				12'd2182	: data2 <= weights[2183];
				12'd2183	: data2 <= weights[2184];
				12'd2184	: data2 <= weights[2185];
				12'd2185	: data2 <= weights[2186];
				12'd2186	: data2 <= weights[2187];
				12'd2187	: data2 <= weights[2188];
				12'd2188	: data2 <= weights[2189];
				12'd2189	: data2 <= weights[2190];
				12'd2190	: data2 <= weights[2191];
				12'd2191	: data2 <= weights[2192];
				12'd2192	: data2 <= weights[2193];
				12'd2193	: data2 <= weights[2194];
				12'd2194	: data2 <= weights[2195];
				12'd2195	: data2 <= weights[2196];
				12'd2196	: data2 <= weights[2197];
				12'd2197	: data2 <= weights[2198];
				12'd2198	: data2 <= weights[2199];
				12'd2199	: data2 <= weights[2200];
				12'd2200	: data2 <= weights[2201];
				12'd2201	: data2 <= weights[2202];
				12'd2202	: data2 <= weights[2203];
				12'd2203	: data2 <= weights[2204];
				12'd2204	: data2 <= weights[2205];
				12'd2205	: data2 <= weights[2206];
				12'd2206	: data2 <= weights[2207];
				12'd2207	: data2 <= weights[2208];
				12'd2208	: data2 <= weights[2209];
				12'd2209	: data2 <= weights[2210];
				12'd2210	: data2 <= weights[2211];
				12'd2211	: data2 <= weights[2212];
				12'd2212	: data2 <= weights[2213];
				12'd2213	: data2 <= weights[2214];
				12'd2214	: data2 <= weights[2215];
				12'd2215	: data2 <= weights[2216];
				12'd2216	: data2 <= weights[2217];
				12'd2217	: data2 <= weights[2218];
				12'd2218	: data2 <= weights[2219];
				12'd2219	: data2 <= weights[2220];
				12'd2220	: data2 <= weights[2221];
				12'd2221	: data2 <= weights[2222];
				12'd2222	: data2 <= weights[2223];
				12'd2223	: data2 <= weights[2224];
				12'd2224	: data2 <= weights[2225];
				12'd2225	: data2 <= weights[2226];
				12'd2226	: data2 <= weights[2227];
				12'd2227	: data2 <= weights[2228];
				12'd2228	: data2 <= weights[2229];
				12'd2229	: data2 <= weights[2230];
				12'd2230	: data2 <= weights[2231];
				12'd2231	: data2 <= weights[2232];
				12'd2232	: data2 <= weights[2233];
				12'd2233	: data2 <= weights[2234];
				12'd2234	: data2 <= weights[2235];
				12'd2235	: data2 <= weights[2236];
				12'd2236	: data2 <= weights[2237];
				12'd2237	: data2 <= weights[2238];
				12'd2238	: data2 <= weights[2239];
				12'd2239	: data2 <= weights[2240];
				12'd2240	: data2 <= weights[2241];
				12'd2241	: data2 <= weights[2242];
				12'd2242	: data2 <= weights[2243];
				12'd2243	: data2 <= weights[2244];
				12'd2244	: data2 <= weights[2245];
				12'd2245	: data2 <= weights[2246];
				12'd2246	: data2 <= weights[2247];
				12'd2247	: data2 <= weights[2248];
				12'd2248	: data2 <= weights[2249];
				12'd2249	: data2 <= weights[2250];
				12'd2250	: data2 <= weights[2251];
				12'd2251	: data2 <= weights[2252];
				12'd2252	: data2 <= weights[2253];
				12'd2253	: data2 <= weights[2254];
				12'd2254	: data2 <= weights[2255];
				12'd2255	: data2 <= weights[2256];
				12'd2256	: data2 <= weights[2257];
				12'd2257	: data2 <= weights[2258];
				12'd2258	: data2 <= weights[2259];
				12'd2259	: data2 <= weights[2260];
				12'd2260	: data2 <= weights[2261];
				12'd2261	: data2 <= weights[2262];
				12'd2262	: data2 <= weights[2263];
				12'd2263	: data2 <= weights[2264];
				12'd2264	: data2 <= weights[2265];
				12'd2265	: data2 <= weights[2266];
				12'd2266	: data2 <= weights[2267];
				12'd2267	: data2 <= weights[2268];
				12'd2268	: data2 <= weights[2269];
				12'd2269	: data2 <= weights[2270];
				12'd2270	: data2 <= weights[2271];
				12'd2271	: data2 <= weights[2272];
				12'd2272	: data2 <= weights[2273];
				12'd2273	: data2 <= weights[2274];
				12'd2274	: data2 <= weights[2275];
				12'd2275	: data2 <= weights[2276];
				12'd2276	: data2 <= weights[2277];
				12'd2277	: data2 <= weights[2278];
				12'd2278	: data2 <= weights[2279];
				12'd2279	: data2 <= weights[2280];
				12'd2280	: data2 <= weights[2281];
				12'd2281	: data2 <= weights[2282];
				12'd2282	: data2 <= weights[2283];
				12'd2283	: data2 <= weights[2284];
				12'd2284	: data2 <= weights[2285];
				12'd2285	: data2 <= weights[2286];
				12'd2286	: data2 <= weights[2287];
				12'd2287	: data2 <= weights[2288];
				12'd2288	: data2 <= weights[2289];
				12'd2289	: data2 <= weights[2290];
				12'd2290	: data2 <= weights[2291];
				12'd2291	: data2 <= weights[2292];
				12'd2292	: data2 <= weights[2293];
				12'd2293	: data2 <= weights[2294];
				12'd2294	: data2 <= weights[2295];
				12'd2295	: data2 <= weights[2296];
				12'd2296	: data2 <= weights[2297];
				12'd2297	: data2 <= weights[2298];
				12'd2298	: data2 <= weights[2299];
				12'd2299	: data2 <= weights[2300];
				12'd2300	: data2 <= weights[2301];
				12'd2301	: data2 <= weights[2302];
				12'd2302	: data2 <= weights[2303];
				12'd2303	: data2 <= weights[2304];
				12'd2304	: data2 <= weights[2305];
				12'd2305	: data2 <= weights[2306];
				12'd2306	: data2 <= weights[2307];
				12'd2307	: data2 <= weights[2308];
				12'd2308	: data2 <= weights[2309];
				12'd2309	: data2 <= weights[2310];
				12'd2310	: data2 <= weights[2311];
				12'd2311	: data2 <= weights[2312];
				12'd2312	: data2 <= weights[2313];
				12'd2313	: data2 <= weights[2314];
				12'd2314	: data2 <= weights[2315];
				12'd2315	: data2 <= weights[2316];
				12'd2316	: data2 <= weights[2317];
				12'd2317	: data2 <= weights[2318];
				12'd2318	: data2 <= weights[2319];
				12'd2319	: data2 <= weights[2320];
				12'd2320	: data2 <= weights[2321];
				12'd2321	: data2 <= weights[2322];
				12'd2322	: data2 <= weights[2323];
				12'd2323	: data2 <= weights[2324];
				12'd2324	: data2 <= weights[2325];
				12'd2325	: data2 <= weights[2326];
				12'd2326	: data2 <= weights[2327];
				12'd2327	: data2 <= weights[2328];
				12'd2328	: data2 <= weights[2329];
				12'd2329	: data2 <= weights[2330];
				12'd2330	: data2 <= weights[2331];
				12'd2331	: data2 <= weights[2332];
				12'd2332	: data2 <= weights[2333];
				12'd2333	: data2 <= weights[2334];
				12'd2334	: data2 <= weights[2335];
				12'd2335	: data2 <= weights[2336];
				12'd2336	: data2 <= weights[2337];
				12'd2337	: data2 <= weights[2338];
				12'd2338	: data2 <= weights[2339];
				12'd2339	: data2 <= weights[2340];
				12'd2340	: data2 <= weights[2341];
				12'd2341	: data2 <= weights[2342];
				12'd2342	: data2 <= weights[2343];
				12'd2343	: data2 <= weights[2344];
				12'd2344	: data2 <= weights[2345];
				12'd2345	: data2 <= weights[2346];
				12'd2346	: data2 <= weights[2347];
				12'd2347	: data2 <= weights[2348];
				12'd2348	: data2 <= weights[2349];
				12'd2349	: data2 <= weights[2350];
				12'd2350	: data2 <= weights[2351];
				12'd2351	: data2 <= weights[2352];
				12'd2352	: data2 <= weights[2353];
				12'd2353	: data2 <= weights[2354];
				12'd2354	: data2 <= weights[2355];
				12'd2355	: data2 <= weights[2356];
				12'd2356	: data2 <= weights[2357];
				12'd2357	: data2 <= weights[2358];
				12'd2358	: data2 <= weights[2359];
				12'd2359	: data2 <= weights[2360];
				12'd2360	: data2 <= weights[2361];
				12'd2361	: data2 <= weights[2362];
				12'd2362	: data2 <= weights[2363];
				12'd2363	: data2 <= weights[2364];
				12'd2364	: data2 <= weights[2365];
				12'd2365	: data2 <= weights[2366];
				12'd2366	: data2 <= weights[2367];
				12'd2367	: data2 <= weights[2368];
				12'd2368	: data2 <= weights[2369];
				12'd2369	: data2 <= weights[2370];
				12'd2370	: data2 <= weights[2371];
				12'd2371	: data2 <= weights[2372];
				12'd2372	: data2 <= weights[2373];
				12'd2373	: data2 <= weights[2374];
				12'd2374	: data2 <= weights[2375];
				12'd2375	: data2 <= weights[2376];
				12'd2376	: data2 <= weights[2377];
				12'd2377	: data2 <= weights[2378];
				12'd2378	: data2 <= weights[2379];
				12'd2379	: data2 <= weights[2380];
				12'd2380	: data2 <= weights[2381];
				12'd2381	: data2 <= weights[2382];
				12'd2382	: data2 <= weights[2383];
				12'd2383	: data2 <= weights[2384];
				12'd2384	: data2 <= weights[2385];
				12'd2385	: data2 <= weights[2386];
				12'd2386	: data2 <= weights[2387];
				12'd2387	: data2 <= weights[2388];
				12'd2388	: data2 <= weights[2389];
				12'd2389	: data2 <= weights[2390];
				12'd2390	: data2 <= weights[2391];
				12'd2391	: data2 <= weights[2392];
				12'd2392	: data2 <= weights[2393];
				12'd2393	: data2 <= weights[2394];
				12'd2394	: data2 <= weights[2395];
				12'd2395	: data2 <= weights[2396];
				12'd2396	: data2 <= weights[2397];
				12'd2397	: data2 <= weights[2398];
				12'd2398	: data2 <= weights[2399];
				12'd2399	: data2 <= weights[2400];
				12'd2400	: data2 <= weights[2401];
				12'd2401	: data2 <= weights[2402];
				12'd2402	: data2 <= weights[2403];
				12'd2403	: data2 <= weights[2404];
				12'd2404	: data2 <= weights[2405];
				12'd2405	: data2 <= weights[2406];
				12'd2406	: data2 <= weights[2407];
				12'd2407	: data2 <= weights[2408];
				12'd2408	: data2 <= weights[2409];
				12'd2409	: data2 <= weights[2410];
				12'd2410	: data2 <= weights[2411];
				12'd2411	: data2 <= weights[2412];
				12'd2412	: data2 <= weights[2413];
				12'd2413	: data2 <= weights[2414];
				12'd2414	: data2 <= weights[2415];
				12'd2415	: data2 <= weights[2416];
				12'd2416	: data2 <= weights[2417];
				12'd2417	: data2 <= weights[2418];
				12'd2418	: data2 <= weights[2419];
				12'd2419	: data2 <= weights[2420];
				12'd2420	: data2 <= weights[2421];
				12'd2421	: data2 <= weights[2422];
				12'd2422	: data2 <= weights[2423];
				12'd2423	: data2 <= weights[2424];
				12'd2424	: data2 <= weights[2425];
				12'd2425	: data2 <= weights[2426];
				12'd2426	: data2 <= weights[2427];
				12'd2427	: data2 <= weights[2428];
				12'd2428	: data2 <= weights[2429];
				12'd2429	: data2 <= weights[2430];
				12'd2430	: data2 <= weights[2431];
				12'd2431	: data2 <= weights[2432];
				12'd2432	: data2 <= weights[2433];
				12'd2433	: data2 <= weights[2434];
				12'd2434	: data2 <= weights[2435];
				12'd2435	: data2 <= weights[2436];
				12'd2436	: data2 <= weights[2437];
				12'd2437	: data2 <= weights[2438];
				12'd2438	: data2 <= weights[2439];
				12'd2439	: data2 <= weights[2440];
				12'd2440	: data2 <= weights[2441];
				12'd2441	: data2 <= weights[2442];
				12'd2442	: data2 <= weights[2443];
				12'd2443	: data2 <= weights[2444];
				12'd2444	: data2 <= weights[2445];
				12'd2445	: data2 <= weights[2446];
				12'd2446	: data2 <= weights[2447];
				12'd2447	: data2 <= weights[2448];
				12'd2448	: data2 <= weights[2449];
				12'd2449	: data2 <= weights[2450];
				12'd2450	: data2 <= weights[2451];
				12'd2451	: data2 <= weights[2452];
				12'd2452	: data2 <= weights[2453];
				12'd2453	: data2 <= weights[2454];
				12'd2454	: data2 <= weights[2455];
				12'd2455	: data2 <= weights[2456];
				12'd2456	: data2 <= weights[2457];
				12'd2457	: data2 <= weights[2458];
				12'd2458	: data2 <= weights[2459];
				12'd2459	: data2 <= weights[2460];
				12'd2460	: data2 <= weights[2461];
				12'd2461	: data2 <= weights[2462];
				12'd2462	: data2 <= weights[2463];
				12'd2463	: data2 <= weights[2464];
				12'd2464	: data2 <= weights[2465];
				12'd2465	: data2 <= weights[2466];
				12'd2466	: data2 <= weights[2467];
				12'd2467	: data2 <= weights[2468];
				12'd2468	: data2 <= weights[2469];
				12'd2469	: data2 <= weights[2470];
				12'd2470	: data2 <= weights[2471];
				12'd2471	: data2 <= weights[2472];
				12'd2472	: data2 <= weights[2473];
				12'd2473	: data2 <= weights[2474];
				12'd2474	: data2 <= weights[2475];
				12'd2475	: data2 <= weights[2476];
				12'd2476	: data2 <= weights[2477];
				12'd2477	: data2 <= weights[2478];
				12'd2478	: data2 <= weights[2479];
				12'd2479	: data2 <= weights[2480];
				12'd2480	: data2 <= weights[2481];
				12'd2481	: data2 <= weights[2482];
				12'd2482	: data2 <= weights[2483];
				12'd2483	: data2 <= weights[2484];
				12'd2484	: data2 <= weights[2485];
				12'd2485	: data2 <= weights[2486];
				12'd2486	: data2 <= weights[2487];
				12'd2487	: data2 <= weights[2488];
				12'd2488	: data2 <= weights[2489];
				12'd2489	: data2 <= weights[2490];
				12'd2490	: data2 <= weights[2491];
				12'd2491	: data2 <= weights[2492];
				12'd2492	: data2 <= weights[2493];
				12'd2493	: data2 <= weights[2494];
				12'd2494	: data2 <= weights[2495];
				12'd2495	: data2 <= weights[2496];
				12'd2496	: data2 <= weights[2497];
				12'd2497	: data2 <= weights[2498];
				12'd2498	: data2 <= weights[2499];
				12'd2499	: data2 <= weights[2500];
				12'd2500	: data2 <= weights[2501];
				12'd2501	: data2 <= weights[2502];
				12'd2502	: data2 <= weights[2503];
				12'd2503	: data2 <= weights[2504];
				12'd2504	: data2 <= weights[2505];
				12'd2505	: data2 <= weights[2506];
				12'd2506	: data2 <= weights[2507];
				12'd2507	: data2 <= weights[2508];
				12'd2508	: data2 <= weights[2509];
				12'd2509	: data2 <= weights[2510];
				12'd2510	: data2 <= weights[2511];
				12'd2511	: data2 <= weights[2512];
				12'd2512	: data2 <= weights[2513];
				12'd2513	: data2 <= weights[2514];
				12'd2514	: data2 <= weights[2515];
				12'd2515	: data2 <= weights[2516];
				12'd2516	: data2 <= weights[2517];
				12'd2517	: data2 <= weights[2518];
				12'd2518	: data2 <= weights[2519];
				12'd2519	: data2 <= weights[2520];
				12'd2520	: data2 <= weights[2521];
				12'd2521	: data2 <= weights[2522];
				12'd2522	: data2 <= weights[2523];
				12'd2523	: data2 <= weights[2524];
				12'd2524	: data2 <= weights[2525];
				12'd2525	: data2 <= weights[2526];
				12'd2526	: data2 <= weights[2527];
				12'd2527	: data2 <= weights[2528];
				12'd2528	: data2 <= weights[2529];
				12'd2529	: data2 <= weights[2530];
				12'd2530	: data2 <= weights[2531];
				12'd2531	: data2 <= weights[2532];
				12'd2532	: data2 <= weights[2533];
				12'd2533	: data2 <= weights[2534];
				12'd2534	: data2 <= weights[2535];
				12'd2535	: data2 <= weights[2536];
				12'd2536	: data2 <= weights[2537];
				12'd2537	: data2 <= weights[2538];
				12'd2538	: data2 <= weights[2539];
				12'd2539	: data2 <= weights[2540];
				12'd2540	: data2 <= weights[2541];
				12'd2541	: data2 <= weights[2542];
				12'd2542	: data2 <= weights[2543];
				12'd2543	: data2 <= weights[2544];
				12'd2544	: data2 <= weights[2545];
				12'd2545	: data2 <= weights[2546];
				12'd2546	: data2 <= weights[2547];
				12'd2547	: data2 <= weights[2548];
				12'd2548	: data2 <= weights[2549];
				12'd2549	: data2 <= weights[2550];
				12'd2550	: data2 <= weights[2551];
				12'd2551	: data2 <= weights[2552];
				12'd2552	: data2 <= weights[2553];
				12'd2553	: data2 <= weights[2554];
				12'd2554	: data2 <= weights[2555];
				12'd2555	: data2 <= weights[2556];
				12'd2556	: data2 <= weights[2557];
				12'd2557	: data2 <= weights[2558];
				12'd2558	: data2 <= weights[2559];
				12'd2559	: data2 <= weights[2560];
				12'd2560	: data2 <= weights[2561];
				12'd2561	: data2 <= weights[2562];
				12'd2562	: data2 <= weights[2563];
				12'd2563	: data2 <= weights[2564];
				12'd2564	: data2 <= weights[2565];
				12'd2565	: data2 <= weights[2566];
				12'd2566	: data2 <= weights[2567];
				12'd2567	: data2 <= weights[2568];
				12'd2568	: data2 <= weights[2569];
				12'd2569	: data2 <= weights[2570];
				12'd2570	: data2 <= weights[2571];
				12'd2571	: data2 <= weights[2572];
				12'd2572	: data2 <= weights[2573];
				12'd2573	: data2 <= weights[2574];
				12'd2574	: data2 <= weights[2575];
				12'd2575	: data2 <= weights[2576];
				12'd2576	: data2 <= weights[2577];
				12'd2577	: data2 <= weights[2578];
				12'd2578	: data2 <= weights[2579];
				12'd2579	: data2 <= weights[2580];
				12'd2580	: data2 <= weights[2581];
				12'd2581	: data2 <= weights[2582];
				12'd2582	: data2 <= weights[2583];
				12'd2583	: data2 <= weights[2584];
				12'd2584	: data2 <= weights[2585];
				12'd2585	: data2 <= weights[2586];
				12'd2586	: data2 <= weights[2587];
				12'd2587	: data2 <= weights[2588];
				12'd2588	: data2 <= weights[2589];
				12'd2589	: data2 <= weights[2590];
				12'd2590	: data2 <= weights[2591];
				12'd2591	: data2 <= weights[2592];
				12'd2592	: data2 <= weights[2593];
				12'd2593	: data2 <= weights[2594];
				12'd2594	: data2 <= weights[2595];
				12'd2595	: data2 <= weights[2596];
				12'd2596	: data2 <= weights[2597];
				12'd2597	: data2 <= weights[2598];
				12'd2598	: data2 <= weights[2599];
				12'd2599	: data2 <= weights[2600];
				12'd2600	: data2 <= weights[2601];
				12'd2601	: data2 <= weights[2602];
				12'd2602	: data2 <= weights[2603];
				12'd2603	: data2 <= weights[2604];
				12'd2604	: data2 <= weights[2605];
				12'd2605	: data2 <= weights[2606];
				12'd2606	: data2 <= weights[2607];
				12'd2607	: data2 <= weights[2608];
				12'd2608	: data2 <= weights[2609];
				12'd2609	: data2 <= weights[2610];
				12'd2610	: data2 <= weights[2611];
				12'd2611	: data2 <= weights[2612];
				12'd2612	: data2 <= weights[2613];
				12'd2613	: data2 <= weights[2614];
				12'd2614	: data2 <= weights[2615];
				12'd2615	: data2 <= weights[2616];
				12'd2616	: data2 <= weights[2617];
				12'd2617	: data2 <= weights[2618];
				12'd2618	: data2 <= weights[2619];
				12'd2619	: data2 <= weights[2620];
				12'd2620	: data2 <= weights[2621];
				12'd2621	: data2 <= weights[2622];
				12'd2622	: data2 <= weights[2623];
				12'd2623	: data2 <= weights[2624];
				12'd2624	: data2 <= weights[2625];
				12'd2625	: data2 <= weights[2626];
				12'd2626	: data2 <= weights[2627];
				12'd2627	: data2 <= weights[2628];
				12'd2628	: data2 <= weights[2629];
				12'd2629	: data2 <= weights[2630];
				12'd2630	: data2 <= weights[2631];
				12'd2631	: data2 <= weights[2632];
				12'd2632	: data2 <= weights[2633];
				12'd2633	: data2 <= weights[2634];
				12'd2634	: data2 <= weights[2635];
				12'd2635	: data2 <= weights[2636];
				12'd2636	: data2 <= weights[2637];
				12'd2637	: data2 <= weights[2638];
				12'd2638	: data2 <= weights[2639];
				12'd2639	: data2 <= weights[2640];
				12'd2640	: data2 <= weights[2641];
				12'd2641	: data2 <= weights[2642];
				12'd2642	: data2 <= weights[2643];
				12'd2643	: data2 <= weights[2644];
				12'd2644	: data2 <= weights[2645];
				12'd2645	: data2 <= weights[2646];
				12'd2646	: data2 <= weights[2647];
				12'd2647	: data2 <= weights[2648];
				12'd2648	: data2 <= weights[2649];
				12'd2649	: data2 <= weights[2650];
				12'd2650	: data2 <= weights[2651];
				12'd2651	: data2 <= weights[2652];
				12'd2652	: data2 <= weights[2653];
				12'd2653	: data2 <= weights[2654];
				12'd2654	: data2 <= weights[2655];
				12'd2655	: data2 <= weights[2656];
				12'd2656	: data2 <= weights[2657];
				12'd2657	: data2 <= weights[2658];
				12'd2658	: data2 <= weights[2659];
				12'd2659	: data2 <= weights[2660];
				12'd2660	: data2 <= weights[2661];
				12'd2661	: data2 <= weights[2662];
				12'd2662	: data2 <= weights[2663];
				12'd2663	: data2 <= weights[2664];
				12'd2664	: data2 <= weights[2665];
				12'd2665	: data2 <= weights[2666];
				12'd2666	: data2 <= weights[2667];
				12'd2667	: data2 <= weights[2668];
				12'd2668	: data2 <= weights[2669];
				12'd2669	: data2 <= weights[2670];
				12'd2670	: data2 <= weights[2671];
				12'd2671	: data2 <= weights[2672];
				12'd2672	: data2 <= weights[2673];
				12'd2673	: data2 <= weights[2674];
				12'd2674	: data2 <= weights[2675];
				12'd2675	: data2 <= weights[2676];
				12'd2676	: data2 <= weights[2677];
				12'd2677	: data2 <= weights[2678];
				12'd2678	: data2 <= weights[2679];
				12'd2679	: data2 <= weights[2680];
				12'd2680	: data2 <= weights[2681];
				12'd2681	: data2 <= weights[2682];
				12'd2682	: data2 <= weights[2683];
				12'd2683	: data2 <= weights[2684];
				12'd2684	: data2 <= weights[2685];
				12'd2685	: data2 <= weights[2686];
				12'd2686	: data2 <= weights[2687];
				12'd2687	: data2 <= weights[2688];
				12'd2688	: data2 <= weights[2689];
				12'd2689	: data2 <= weights[2690];
				12'd2690	: data2 <= weights[2691];
				12'd2691	: data2 <= weights[2692];
				12'd2692	: data2 <= weights[2693];
				12'd2693	: data2 <= weights[2694];
				12'd2694	: data2 <= weights[2695];
				12'd2695	: data2 <= weights[2696];
				12'd2696	: data2 <= weights[2697];
				12'd2697	: data2 <= weights[2698];
				12'd2698	: data2 <= weights[2699];
				12'd2699	: data2 <= weights[2700];
				12'd2700	: data2 <= weights[2701];
				12'd2701	: data2 <= weights[2702];
				12'd2702	: data2 <= weights[2703];
				12'd2703	: data2 <= weights[2704];
				12'd2704	: data2 <= weights[2705];
				12'd2705	: data2 <= weights[2706];
				12'd2706	: data2 <= weights[2707];
				12'd2707	: data2 <= weights[2708];
				12'd2708	: data2 <= weights[2709];
				12'd2709	: data2 <= weights[2710];
				12'd2710	: data2 <= weights[2711];
				12'd2711	: data2 <= weights[2712];
				12'd2712	: data2 <= weights[2713];
				12'd2713	: data2 <= weights[2714];
				12'd2714	: data2 <= weights[2715];
				12'd2715	: data2 <= weights[2716];
				12'd2716	: data2 <= weights[2717];
				12'd2717	: data2 <= weights[2718];
				12'd2718	: data2 <= weights[2719];
				12'd2719	: data2 <= weights[2720];
				12'd2720	: data2 <= weights[2721];
				12'd2721	: data2 <= weights[2722];
				12'd2722	: data2 <= weights[2723];
				12'd2723	: data2 <= weights[2724];
				12'd2724	: data2 <= weights[2725];
				12'd2725	: data2 <= weights[2726];
				12'd2726	: data2 <= weights[2727];
				12'd2727	: data2 <= weights[2728];
				12'd2728	: data2 <= weights[2729];
				12'd2729	: data2 <= weights[2730];
				12'd2730	: data2 <= weights[2731];
				12'd2731	: data2 <= weights[2732];
				12'd2732	: data2 <= weights[2733];
				12'd2733	: data2 <= weights[2734];
				12'd2734	: data2 <= weights[2735];
				12'd2735	: data2 <= weights[2736];
				12'd2736	: data2 <= weights[2737];
				12'd2737	: data2 <= weights[2738];
				12'd2738	: data2 <= weights[2739];
				12'd2739	: data2 <= weights[2740];
				12'd2740	: data2 <= weights[2741];
				12'd2741	: data2 <= weights[2742];
				12'd2742	: data2 <= weights[2743];
				12'd2743	: data2 <= weights[2744];
				12'd2744	: data2 <= weights[2745];
				12'd2745	: data2 <= weights[2746];
				12'd2746	: data2 <= weights[2747];
				12'd2747	: data2 <= weights[2748];
				12'd2748	: data2 <= weights[2749];
				12'd2749	: data2 <= weights[2750];
				12'd2750	: data2 <= weights[2751];
				12'd2751	: data2 <= weights[2752];
				12'd2752	: data2 <= weights[2753];
				12'd2753	: data2 <= weights[2754];
				12'd2754	: data2 <= weights[2755];
				12'd2755	: data2 <= weights[2756];
				12'd2756	: data2 <= weights[2757];
				12'd2757	: data2 <= weights[2758];
				12'd2758	: data2 <= weights[2759];
				12'd2759	: data2 <= weights[2760];
				12'd2760	: data2 <= weights[2761];
				12'd2761	: data2 <= weights[2762];
				12'd2762	: data2 <= weights[2763];
				12'd2763	: data2 <= weights[2764];
				12'd2764	: data2 <= weights[2765];
				12'd2765	: data2 <= weights[2766];
				12'd2766	: data2 <= weights[2767];
				12'd2767	: data2 <= weights[2768];
				12'd2768	: data2 <= weights[2769];
				12'd2769	: data2 <= weights[2770];
				12'd2770	: data2 <= weights[2771];
				12'd2771	: data2 <= weights[2772];
				12'd2772	: data2 <= weights[2773];
				12'd2773	: data2 <= weights[2774];
				12'd2774	: data2 <= weights[2775];
				12'd2775	: data2 <= weights[2776];
				12'd2776	: data2 <= weights[2777];
				12'd2777	: data2 <= weights[2778];
				12'd2778	: data2 <= weights[2779];
				12'd2779	: data2 <= weights[2780];
				12'd2780	: data2 <= weights[2781];
				12'd2781	: data2 <= weights[2782];
				12'd2782	: data2 <= weights[2783];
				12'd2783	: data2 <= weights[2784];
				12'd2784	: data2 <= weights[2785];
				12'd2785	: data2 <= weights[2786];
				12'd2786	: data2 <= weights[2787];
				12'd2787	: data2 <= weights[2788];
				12'd2788	: data2 <= weights[2789];
				12'd2789	: data2 <= weights[2790];
				12'd2790	: data2 <= weights[2791];
				12'd2791	: data2 <= weights[2792];
				12'd2792	: data2 <= weights[2793];
				12'd2793	: data2 <= weights[2794];
				12'd2794	: data2 <= weights[2795];
				12'd2795	: data2 <= weights[2796];
				12'd2796	: data2 <= weights[2797];
				12'd2797	: data2 <= weights[2798];
				12'd2798	: data2 <= weights[2799];
				12'd2799	: data2 <= weights[2800];
				12'd2800	: data2 <= weights[2801];
				12'd2801	: data2 <= weights[2802];
				12'd2802	: data2 <= weights[2803];
				12'd2803	: data2 <= weights[2804];
				12'd2804	: data2 <= weights[2805];
				12'd2805	: data2 <= weights[2806];
				12'd2806	: data2 <= weights[2807];
				12'd2807	: data2 <= weights[2808];
				12'd2808	: data2 <= weights[2809];
				12'd2809	: data2 <= weights[2810];
				12'd2810	: data2 <= weights[2811];
				12'd2811	: data2 <= weights[2812];
				12'd2812	: data2 <= weights[2813];
				12'd2813	: data2 <= weights[2814];
				12'd2814	: data2 <= weights[2815];
				12'd2815	: data2 <= weights[2816];
				12'd2816	: data2 <= weights[2817];
				12'd2817	: data2 <= weights[2818];
				12'd2818	: data2 <= weights[2819];
				12'd2819	: data2 <= weights[2820];
				12'd2820	: data2 <= weights[2821];
				12'd2821	: data2 <= weights[2822];
				12'd2822	: data2 <= weights[2823];
				12'd2823	: data2 <= weights[2824];
				12'd2824	: data2 <= weights[2825];
				12'd2825	: data2 <= weights[2826];
				12'd2826	: data2 <= weights[2827];
				12'd2827	: data2 <= weights[2828];
				12'd2828	: data2 <= weights[2829];
				12'd2829	: data2 <= weights[2830];
				12'd2830	: data2 <= weights[2831];
				12'd2831	: data2 <= weights[2832];
				12'd2832	: data2 <= weights[2833];
				12'd2833	: data2 <= weights[2834];
				12'd2834	: data2 <= weights[2835];
				12'd2835	: data2 <= weights[2836];
				12'd2836	: data2 <= weights[2837];
				12'd2837	: data2 <= weights[2838];
				12'd2838	: data2 <= weights[2839];
				12'd2839	: data2 <= weights[2840];
				12'd2840	: data2 <= weights[2841];
				12'd2841	: data2 <= weights[2842];
				12'd2842	: data2 <= weights[2843];
				12'd2843	: data2 <= weights[2844];
				12'd2844	: data2 <= weights[2845];
				12'd2845	: data2 <= weights[2846];
				12'd2846	: data2 <= weights[2847];
				12'd2847	: data2 <= weights[2848];
				12'd2848	: data2 <= weights[2849];
				12'd2849	: data2 <= weights[2850];
				12'd2850	: data2 <= weights[2851];
				12'd2851	: data2 <= weights[2852];
				12'd2852	: data2 <= weights[2853];
				12'd2853	: data2 <= weights[2854];
				12'd2854	: data2 <= weights[2855];
				12'd2855	: data2 <= weights[2856];
				12'd2856	: data2 <= weights[2857];
				12'd2857	: data2 <= weights[2858];
				12'd2858	: data2 <= weights[2859];
				12'd2859	: data2 <= weights[2860];
				12'd2860	: data2 <= weights[2861];
				12'd2861	: data2 <= weights[2862];
				12'd2862	: data2 <= weights[2863];
				12'd2863	: data2 <= weights[2864];
				12'd2864	: data2 <= weights[2865];
				12'd2865	: data2 <= weights[2866];
				12'd2866	: data2 <= weights[2867];
				12'd2867	: data2 <= weights[2868];
				12'd2868	: data2 <= weights[2869];
				12'd2869	: data2 <= weights[2870];
				12'd2870	: data2 <= weights[2871];
				12'd2871	: data2 <= weights[2872];
				12'd2872	: data2 <= weights[2873];
				12'd2873	: data2 <= weights[2874];
				12'd2874	: data2 <= weights[2875];
				12'd2875	: data2 <= weights[2876];
				12'd2876	: data2 <= weights[2877];
				12'd2877	: data2 <= weights[2878];
				12'd2878	: data2 <= weights[2879];
				12'd2879	: data2 <= weights[2880];
				12'd2880	: data2 <= weights[2881];
				12'd2881	: data2 <= weights[2882];
				12'd2882	: data2 <= weights[2883];
				12'd2883	: data2 <= weights[2884];
				12'd2884	: data2 <= weights[2885];
				12'd2885	: data2 <= weights[2886];
				12'd2886	: data2 <= weights[2887];
				12'd2887	: data2 <= weights[2888];
				12'd2888	: data2 <= weights[2889];
				12'd2889	: data2 <= weights[2890];
				12'd2890	: data2 <= weights[2891];
				12'd2891	: data2 <= weights[2892];
				12'd2892	: data2 <= weights[2893];
				12'd2893	: data2 <= weights[2894];
				12'd2894	: data2 <= weights[2895];
				12'd2895	: data2 <= weights[2896];
				12'd2896	: data2 <= weights[2897];
				12'd2897	: data2 <= weights[2898];
				12'd2898	: data2 <= weights[2899];
				12'd2899	: data2 <= weights[2900];
				12'd2900	: data2 <= weights[2901];
				12'd2901	: data2 <= weights[2902];
				12'd2902	: data2 <= weights[2903];
				12'd2903	: data2 <= weights[2904];
				12'd2904	: data2 <= weights[2905];
				12'd2905	: data2 <= weights[2906];
				12'd2906	: data2 <= weights[2907];
				12'd2907	: data2 <= weights[2908];
				12'd2908	: data2 <= weights[2909];
				12'd2909	: data2 <= weights[2910];
				12'd2910	: data2 <= weights[2911];
				12'd2911	: data2 <= weights[2912];
				12'd2912	: data2 <= weights[2913];
				12'd2913	: data2 <= weights[2914];
				12'd2914	: data2 <= weights[2915];
				12'd2915	: data2 <= weights[2916];
				12'd2916	: data2 <= weights[2917];
				12'd2917	: data2 <= weights[2918];
				12'd2918	: data2 <= weights[2919];
				12'd2919	: data2 <= weights[2920];
				12'd2920	: data2 <= weights[2921];
				12'd2921	: data2 <= weights[2922];
				12'd2922	: data2 <= weights[2923];
				12'd2923	: data2 <= weights[2924];
				12'd2924	: data2 <= weights[2925];
				12'd2925	: data2 <= weights[2926];
				12'd2926	: data2 <= weights[2927];
				12'd2927	: data2 <= weights[2928];
				12'd2928	: data2 <= weights[2929];
				12'd2929	: data2 <= weights[2930];
				12'd2930	: data2 <= weights[2931];
				12'd2931	: data2 <= weights[2932];
				12'd2932	: data2 <= weights[2933];
				12'd2933	: data2 <= weights[2934];
				12'd2934	: data2 <= weights[2935];
				12'd2935	: data2 <= weights[2936];
				12'd2936	: data2 <= weights[2937];
				12'd2937	: data2 <= weights[2938];
				12'd2938	: data2 <= weights[2939];
				12'd2939	: data2 <= weights[2940];
				12'd2940	: data2 <= weights[2941];
				12'd2941	: data2 <= weights[2942];
				12'd2942	: data2 <= weights[2943];
				12'd2943	: data2 <= weights[2944];
				12'd2944	: data2 <= weights[2945];
				12'd2945	: data2 <= weights[2946];
				12'd2946	: data2 <= weights[2947];
				12'd2947	: data2 <= weights[2948];
				12'd2948	: data2 <= weights[2949];
				12'd2949	: data2 <= weights[2950];
				12'd2950	: data2 <= weights[2951];
				12'd2951	: data2 <= weights[2952];
				12'd2952	: data2 <= weights[2953];
				12'd2953	: data2 <= weights[2954];
				12'd2954	: data2 <= weights[2955];
				12'd2955	: data2 <= weights[2956];
				12'd2956	: data2 <= weights[2957];
				12'd2957	: data2 <= weights[2958];
				12'd2958	: data2 <= weights[2959];
				12'd2959	: data2 <= weights[2960];
				12'd2960	: data2 <= weights[2961];
				12'd2961	: data2 <= weights[2962];
				12'd2962	: data2 <= weights[2963];
				12'd2963	: data2 <= weights[2964];
				12'd2964	: data2 <= weights[2965];
				12'd2965	: data2 <= weights[2966];
				12'd2966	: data2 <= weights[2967];
				12'd2967	: data2 <= weights[2968];
				12'd2968	: data2 <= weights[2969];
				12'd2969	: data2 <= weights[2970];
				12'd2970	: data2 <= weights[2971];
				12'd2971	: data2 <= weights[2972];
				12'd2972	: data2 <= weights[2973];
				12'd2973	: data2 <= weights[2974];
				12'd2974	: data2 <= weights[2975];
				12'd2975	: data2 <= weights[2976];
				12'd2976	: data2 <= weights[2977];
				12'd2977	: data2 <= weights[2978];
				12'd2978	: data2 <= weights[2979];
				12'd2979	: data2 <= weights[2980];
				12'd2980	: data2 <= weights[2981];
				12'd2981	: data2 <= weights[2982];
				12'd2982	: data2 <= weights[2983];
				12'd2983	: data2 <= weights[2984];
				12'd2984	: data2 <= weights[2985];
				12'd2985	: data2 <= weights[2986];
				12'd2986	: data2 <= weights[2987];
				12'd2987	: data2 <= weights[2988];
				12'd2988	: data2 <= weights[2989];
				12'd2989	: data2 <= weights[2990];
				12'd2990	: data2 <= weights[2991];
				12'd2991	: data2 <= weights[2992];
				12'd2992	: data2 <= weights[2993];
				12'd2993	: data2 <= weights[2994];
				12'd2994	: data2 <= weights[2995];
				12'd2995	: data2 <= weights[2996];
				12'd2996	: data2 <= weights[2997];
				12'd2997	: data2 <= weights[2998];
				12'd2998	: data2 <= weights[2999];
				12'd2999	: data2 <= weights[3000];
				12'd3000	: data2 <= weights[3001];
				12'd3001	: data2 <= weights[3002];
				12'd3002	: data2 <= weights[3003];
				12'd3003	: data2 <= weights[3004];
				12'd3004	: data2 <= weights[3005];
				12'd3005	: data2 <= weights[3006];
				12'd3006	: data2 <= weights[3007];
				12'd3007	: data2 <= weights[3008];
				12'd3008	: data2 <= weights[3009];
				12'd3009	: data2 <= weights[3010];
				12'd3010	: data2 <= weights[3011];
				12'd3011	: data2 <= weights[3012];
				12'd3012	: data2 <= weights[3013];
				12'd3013	: data2 <= weights[3014];
				12'd3014	: data2 <= weights[3015];
				12'd3015	: data2 <= weights[3016];
				12'd3016	: data2 <= weights[3017];
				12'd3017	: data2 <= weights[3018];
				12'd3018	: data2 <= weights[3019];
				12'd3019	: data2 <= weights[3020];
				12'd3020	: data2 <= weights[3021];
				12'd3021	: data2 <= weights[3022];
				12'd3022	: data2 <= weights[3023];
				12'd3023	: data2 <= weights[3024];
				12'd3024	: data2 <= weights[3025];
				12'd3025	: data2 <= weights[3026];
				12'd3026	: data2 <= weights[3027];
				12'd3027	: data2 <= weights[3028];
				12'd3028	: data2 <= weights[3029];
				12'd3029	: data2 <= weights[3030];
				12'd3030	: data2 <= weights[3031];
				12'd3031	: data2 <= weights[3032];
				12'd3032	: data2 <= weights[3033];
				12'd3033	: data2 <= weights[3034];
				12'd3034	: data2 <= weights[3035];
				12'd3035	: data2 <= weights[3036];
				12'd3036	: data2 <= weights[3037];
				12'd3037	: data2 <= weights[3038];
				12'd3038	: data2 <= weights[3039];
				12'd3039	: data2 <= weights[3040];
				12'd3040	: data2 <= weights[3041];
				12'd3041	: data2 <= weights[3042];
				12'd3042	: data2 <= weights[3043];
				12'd3043	: data2 <= weights[3044];
				12'd3044	: data2 <= weights[3045];
				12'd3045	: data2 <= weights[3046];
				12'd3046	: data2 <= weights[3047];
				12'd3047	: data2 <= weights[3048];
				12'd3048	: data2 <= weights[3049];
				12'd3049	: data2 <= weights[3050];
				12'd3050	: data2 <= weights[3051];
				12'd3051	: data2 <= weights[3052];
				12'd3052	: data2 <= weights[3053];
				12'd3053	: data2 <= weights[3054];
				12'd3054	: data2 <= weights[3055];
				12'd3055	: data2 <= weights[3056];
				12'd3056	: data2 <= weights[3057];
				12'd3057	: data2 <= weights[3058];
				12'd3058	: data2 <= weights[3059];
				12'd3059	: data2 <= weights[3060];
				12'd3060	: data2 <= weights[3061];
				12'd3061	: data2 <= weights[3062];
				12'd3062	: data2 <= weights[3063];
				12'd3063	: data2 <= weights[3064];
				12'd3064	: data2 <= weights[3065];
				12'd3065	: data2 <= weights[3066];
				12'd3066	: data2 <= weights[3067];
				12'd3067	: data2 <= weights[3068];
				12'd3068	: data2 <= weights[3069];
				12'd3069	: data2 <= weights[3070];
				12'd3070	: data2 <= weights[3071];
				12'd3071	: data2 <= weights[3072];
				12'd3072	: data2 <= weights[3073];
				12'd3073	: data2 <= weights[3074];
				12'd3074	: data2 <= weights[3075];
				12'd3075	: data2 <= weights[3076];
				12'd3076	: data2 <= weights[3077];
				12'd3077	: data2 <= weights[3078];
				12'd3078	: data2 <= weights[3079];
				12'd3079	: data2 <= weights[3080];
				12'd3080	: data2 <= weights[3081];
				12'd3081	: data2 <= weights[3082];
				12'd3082	: data2 <= weights[3083];
				12'd3083	: data2 <= weights[3084];
				12'd3084	: data2 <= weights[3085];
				12'd3085	: data2 <= weights[3086];
				12'd3086	: data2 <= weights[3087];
				12'd3087	: data2 <= weights[3088];
				12'd3088	: data2 <= weights[3089];
				12'd3089	: data2 <= weights[3090];
				12'd3090	: data2 <= weights[3091];
				12'd3091	: data2 <= weights[3092];
				12'd3092	: data2 <= weights[3093];
				12'd3093	: data2 <= weights[3094];
				12'd3094	: data2 <= weights[3095];
				12'd3095	: data2 <= weights[3096];
				12'd3096	: data2 <= weights[3097];
				12'd3097	: data2 <= weights[3098];
				12'd3098	: data2 <= weights[3099];
				12'd3099	: data2 <= weights[3100];
				12'd3100	: data2 <= weights[3101];
				12'd3101	: data2 <= weights[3102];
				12'd3102	: data2 <= weights[3103];
				12'd3103	: data2 <= weights[3104];
				12'd3104	: data2 <= weights[3105];
				12'd3105	: data2 <= weights[3106];
				12'd3106	: data2 <= weights[3107];
				12'd3107	: data2 <= weights[3108];
				12'd3108	: data2 <= weights[3109];
				12'd3109	: data2 <= weights[3110];
				12'd3110	: data2 <= weights[3111];
				12'd3111	: data2 <= weights[3112];
				12'd3112	: data2 <= weights[3113];
				12'd3113	: data2 <= weights[3114];
				12'd3114	: data2 <= weights[3115];
				12'd3115	: data2 <= weights[3116];
				12'd3116	: data2 <= weights[3117];
				12'd3117	: data2 <= weights[3118];
				12'd3118	: data2 <= weights[3119];
				12'd3119	: data2 <= weights[3120];
				12'd3120	: data2 <= weights[3121];
				12'd3121	: data2 <= weights[3122];
				12'd3122	: data2 <= weights[3123];
				12'd3123	: data2 <= weights[3124];
				12'd3124	: data2 <= weights[3125];
				12'd3125	: data2 <= weights[3126];
				12'd3126	: data2 <= weights[3127];
				12'd3127	: data2 <= weights[3128];
				12'd3128	: data2 <= weights[3129];
				12'd3129	: data2 <= weights[3130];
				12'd3130	: data2 <= weights[3131];
				12'd3131	: data2 <= weights[3132];
				12'd3132	: data2 <= weights[3133];
				12'd3133	: data2 <= weights[3134];
				12'd3134	: data2 <= weights[3135];
				12'd3135	: data2 <= weights[3136];
				12'd3136	: data2 <= weights[3137];
				12'd3137	: data2 <= weights[3138];
				12'd3138	: data2 <= weights[3139];
				12'd3139	: data2 <= weights[3140];
				12'd3140	: data2 <= weights[3141];
				12'd3141	: data2 <= weights[3142];
				12'd3142	: data2 <= weights[3143];
				12'd3143	: data2 <= weights[3144];
				12'd3144	: data2 <= weights[3145];
				12'd3145	: data2 <= weights[3146];
				12'd3146	: data2 <= weights[3147];
				12'd3147	: data2 <= weights[3148];
				12'd3148	: data2 <= weights[3149];
				12'd3149	: data2 <= weights[3150];
				12'd3150	: data2 <= weights[3151];
				12'd3151	: data2 <= weights[3152];
				12'd3152	: data2 <= weights[3153];
				12'd3153	: data2 <= weights[3154];
				12'd3154	: data2 <= weights[3155];
				12'd3155	: data2 <= weights[3156];
				12'd3156	: data2 <= weights[3157];
				12'd3157	: data2 <= weights[3158];
				12'd3158	: data2 <= weights[3159];
				12'd3159	: data2 <= weights[3160];
				12'd3160	: data2 <= weights[3161];
				12'd3161	: data2 <= weights[3162];
				12'd3162	: data2 <= weights[3163];
				12'd3163	: data2 <= weights[3164];
				12'd3164	: data2 <= weights[3165];
				12'd3165	: data2 <= weights[3166];
				12'd3166	: data2 <= weights[3167];
				12'd3167	: data2 <= weights[3168];
				12'd3168	: data2 <= weights[3169];
				12'd3169	: data2 <= weights[3170];
				12'd3170	: data2 <= weights[3171];
				12'd3171	: data2 <= weights[3172];
				12'd3172	: data2 <= weights[3173];
				12'd3173	: data2 <= weights[3174];
				12'd3174	: data2 <= weights[3175];
				12'd3175	: data2 <= weights[3176];
				12'd3176	: data2 <= weights[3177];
				12'd3177	: data2 <= weights[3178];
				12'd3178	: data2 <= weights[3179];
				12'd3179	: data2 <= weights[3180];
				12'd3180	: data2 <= weights[3181];
				12'd3181	: data2 <= weights[3182];
				12'd3182	: data2 <= weights[3183];
				12'd3183	: data2 <= weights[3184];
				12'd3184	: data2 <= weights[3185];
				12'd3185	: data2 <= weights[3186];
				12'd3186	: data2 <= weights[3187];
				12'd3187	: data2 <= weights[3188];
				12'd3188	: data2 <= weights[3189];
				12'd3189	: data2 <= weights[3190];
				12'd3190	: data2 <= weights[3191];
				12'd3191	: data2 <= weights[3192];
				12'd3192	: data2 <= weights[3193];
				12'd3193	: data2 <= weights[3194];
				12'd3194	: data2 <= weights[3195];
				12'd3195	: data2 <= weights[3196];
				12'd3196	: data2 <= weights[3197];
				12'd3197	: data2 <= weights[3198];
				12'd3198	: data2 <= weights[3199];
				12'd3199	: data2 <= weights[3200];
				12'd3200	: data2 <= weights[3201];
				12'd3201	: data2 <= weights[3202];
				12'd3202	: data2 <= weights[3203];
				12'd3203	: data2 <= weights[3204];
				12'd3204	: data2 <= weights[3205];
				12'd3205	: data2 <= weights[3206];
				12'd3206	: data2 <= weights[3207];
				12'd3207	: data2 <= weights[3208];
				12'd3208	: data2 <= weights[3209];
				12'd3209	: data2 <= weights[3210];
				12'd3210	: data2 <= weights[3211];
				12'd3211	: data2 <= weights[3212];
				12'd3212	: data2 <= weights[3213];
				12'd3213	: data2 <= weights[3214];
				12'd3214	: data2 <= weights[3215];
				12'd3215	: data2 <= weights[3216];
				12'd3216	: data2 <= weights[3217];
				12'd3217	: data2 <= weights[3218];
				12'd3218	: data2 <= weights[3219];
				12'd3219	: data2 <= weights[3220];
				12'd3220	: data2 <= weights[3221];
				12'd3221	: data2 <= weights[3222];
				12'd3222	: data2 <= weights[3223];
				12'd3223	: data2 <= weights[3224];
				12'd3224	: data2 <= weights[3225];
				12'd3225	: data2 <= weights[3226];
				12'd3226	: data2 <= weights[3227];
				12'd3227	: data2 <= weights[3228];
				12'd3228	: data2 <= weights[3229];
				12'd3229	: data2 <= weights[3230];
				12'd3230	: data2 <= weights[3231];
				12'd3231	: data2 <= weights[3232];
				12'd3232	: data2 <= weights[3233];
				12'd3233	: data2 <= weights[3234];
				12'd3234	: data2 <= weights[3235];
				12'd3235	: data2 <= weights[3236];
				12'd3236	: data2 <= weights[3237];
				12'd3237	: data2 <= weights[3238];
				12'd3238	: data2 <= weights[3239];
				12'd3239	: data2 <= weights[3240];
				12'd3240	: data2 <= weights[3241];
				12'd3241	: data2 <= weights[3242];
				12'd3242	: data2 <= weights[3243];
				12'd3243	: data2 <= weights[3244];
				12'd3244	: data2 <= weights[3245];
				12'd3245	: data2 <= weights[3246];
				12'd3246	: data2 <= weights[3247];
				12'd3247	: data2 <= weights[3248];
				12'd3248	: data2 <= weights[3249];
				12'd3249	: data2 <= weights[3250];
				12'd3250	: data2 <= weights[3251];
				12'd3251	: data2 <= weights[3252];
				12'd3252	: data2 <= weights[3253];
				12'd3253	: data2 <= weights[3254];
				12'd3254	: data2 <= weights[3255];
				12'd3255	: data2 <= weights[3256];
				12'd3256	: data2 <= weights[3257];
				12'd3257	: data2 <= weights[3258];
				12'd3258	: data2 <= weights[3259];
				12'd3259	: data2 <= weights[3260];
				12'd3260	: data2 <= weights[3261];
				12'd3261	: data2 <= weights[3262];
				12'd3262	: data2 <= weights[3263];
				12'd3263	: data2 <= weights[3264];
				12'd3264	: data2 <= weights[3265];
				12'd3265	: data2 <= weights[3266];
				12'd3266	: data2 <= weights[3267];
				12'd3267	: data2 <= weights[3268];
				12'd3268	: data2 <= weights[3269];
				12'd3269	: data2 <= weights[3270];
				12'd3270	: data2 <= weights[3271];
				12'd3271	: data2 <= weights[3272];
				12'd3272	: data2 <= weights[3273];
				12'd3273	: data2 <= weights[3274];
				12'd3274	: data2 <= weights[3275];
				12'd3275	: data2 <= weights[3276];
				12'd3276	: data2 <= weights[3277];
				12'd3277	: data2 <= weights[3278];
				12'd3278	: data2 <= weights[3279];
				12'd3279	: data2 <= weights[3280];
				12'd3280	: data2 <= weights[3281];
				12'd3281	: data2 <= weights[3282];
				12'd3282	: data2 <= weights[3283];
				12'd3283	: data2 <= weights[3284];
				12'd3284	: data2 <= weights[3285];
				12'd3285	: data2 <= weights[3286];
				12'd3286	: data2 <= weights[3287];
				12'd3287	: data2 <= weights[3288];
				12'd3288	: data2 <= weights[3289];
				12'd3289	: data2 <= weights[3290];
				12'd3290	: data2 <= weights[3291];
				12'd3291	: data2 <= weights[3292];
				12'd3292	: data2 <= weights[3293];
				12'd3293	: data2 <= weights[3294];
				12'd3294	: data2 <= weights[3295];
				12'd3295	: data2 <= weights[3296];
				12'd3296	: data2 <= weights[3297];
				12'd3297	: data2 <= weights[3298];
				12'd3298	: data2 <= weights[3299];
				12'd3299	: data2 <= weights[3300];
				12'd3300	: data2 <= weights[3301];
				12'd3301	: data2 <= weights[3302];
				12'd3302	: data2 <= weights[3303];
				12'd3303	: data2 <= weights[3304];
				12'd3304	: data2 <= weights[3305];
				12'd3305	: data2 <= weights[3306];
				12'd3306	: data2 <= weights[3307];
				12'd3307	: data2 <= weights[3308];
				12'd3308	: data2 <= weights[3309];
				12'd3309	: data2 <= weights[3310];
				12'd3310	: data2 <= weights[3311];
				12'd3311	: data2 <= weights[3312];
				12'd3312	: data2 <= weights[3313];
				12'd3313	: data2 <= weights[3314];
				12'd3314	: data2 <= weights[3315];
				12'd3315	: data2 <= weights[3316];
				12'd3316	: data2 <= weights[3317];
				12'd3317	: data2 <= weights[3318];
				12'd3318	: data2 <= weights[3319];
				12'd3319	: data2 <= weights[3320];
				12'd3320	: data2 <= weights[3321];
				12'd3321	: data2 <= weights[3322];
				12'd3322	: data2 <= weights[3323];
				12'd3323	: data2 <= weights[3324];
				12'd3324	: data2 <= weights[3325];
				12'd3325	: data2 <= weights[3326];
				12'd3326	: data2 <= weights[3327];
				12'd3327	: data2 <= weights[3328];
				12'd3328	: data2 <= weights[3329];
				12'd3329	: data2 <= weights[3330];
				12'd3330	: data2 <= weights[3331];
				12'd3331	: data2 <= weights[3332];
				12'd3332	: data2 <= weights[3333];
				12'd3333	: data2 <= weights[3334];
				12'd3334	: data2 <= weights[3335];
				12'd3335	: data2 <= weights[3336];
				12'd3336	: data2 <= weights[3337];
				12'd3337	: data2 <= weights[3338];
				12'd3338	: data2 <= weights[3339];
				12'd3339	: data2 <= weights[3340];
				12'd3340	: data2 <= weights[3341];
				12'd3341	: data2 <= weights[3342];
				12'd3342	: data2 <= weights[3343];
				12'd3343	: data2 <= weights[3344];
				12'd3344	: data2 <= weights[3345];
				12'd3345	: data2 <= weights[3346];
				12'd3346	: data2 <= weights[3347];
				12'd3347	: data2 <= weights[3348];
				12'd3348	: data2 <= weights[3349];
				12'd3349	: data2 <= weights[3350];
				12'd3350	: data2 <= weights[3351];
				12'd3351	: data2 <= weights[3352];
				12'd3352	: data2 <= weights[3353];
				12'd3353	: data2 <= weights[3354];
				12'd3354	: data2 <= weights[3355];
				12'd3355	: data2 <= weights[3356];
				12'd3356	: data2 <= weights[3357];
				12'd3357	: data2 <= weights[3358];
				12'd3358	: data2 <= weights[3359];
				12'd3359	: data2 <= weights[3360];
				12'd3360	: data2 <= weights[3361];
				12'd3361	: data2 <= weights[3362];
				12'd3362	: data2 <= weights[3363];
				12'd3363	: data2 <= weights[3364];
				12'd3364	: data2 <= weights[3365];
				12'd3365	: data2 <= weights[3366];
				12'd3366	: data2 <= weights[3367];
				12'd3367	: data2 <= weights[3368];
				12'd3368	: data2 <= weights[3369];
				12'd3369	: data2 <= weights[3370];
				12'd3370	: data2 <= weights[3371];
				12'd3371	: data2 <= weights[3372];
				12'd3372	: data2 <= weights[3373];
				12'd3373	: data2 <= weights[3374];
				12'd3374	: data2 <= weights[3375];
				12'd3375	: data2 <= weights[3376];
				12'd3376	: data2 <= weights[3377];
				12'd3377	: data2 <= weights[3378];
				12'd3378	: data2 <= weights[3379];
				12'd3379	: data2 <= weights[3380];
				12'd3380	: data2 <= weights[3381];
				12'd3381	: data2 <= weights[3382];
				12'd3382	: data2 <= weights[3383];
				12'd3383	: data2 <= weights[3384];
				12'd3384	: data2 <= weights[3385];
				12'd3385	: data2 <= weights[3386];
				12'd3386	: data2 <= weights[3387];
				12'd3387	: data2 <= weights[3388];
				12'd3388	: data2 <= weights[3389];
				12'd3389	: data2 <= weights[3390];
				12'd3390	: data2 <= weights[3391];
				12'd3391	: data2 <= weights[3392];
				12'd3392	: data2 <= weights[3393];
				12'd3393	: data2 <= weights[3394];
				12'd3394	: data2 <= weights[3395];
				12'd3395	: data2 <= weights[3396];
				12'd3396	: data2 <= weights[3397];
				12'd3397	: data2 <= weights[3398];
				12'd3398	: data2 <= weights[3399];
				12'd3399	: data2 <= weights[3400];
				12'd3400	: data2 <= weights[3401];
				12'd3401	: data2 <= weights[3402];
				12'd3402	: data2 <= weights[3403];
				12'd3403	: data2 <= weights[3404];
				12'd3404	: data2 <= weights[3405];
				12'd3405	: data2 <= weights[3406];
				12'd3406	: data2 <= weights[3407];
				12'd3407	: data2 <= weights[3408];
				12'd3408	: data2 <= weights[3409];
				12'd3409	: data2 <= weights[3410];
				12'd3410	: data2 <= weights[3411];
				12'd3411	: data2 <= weights[3412];
				12'd3412	: data2 <= weights[3413];
				12'd3413	: data2 <= weights[3414];
				12'd3414	: data2 <= weights[3415];
				12'd3415	: data2 <= weights[3416];
				12'd3416	: data2 <= weights[3417];
				12'd3417	: data2 <= weights[3418];
				12'd3418	: data2 <= weights[3419];
				12'd3419	: data2 <= weights[3420];
				12'd3420	: data2 <= weights[3421];
				12'd3421	: data2 <= weights[3422];
				12'd3422	: data2 <= weights[3423];
				12'd3423	: data2 <= weights[3424];
				12'd3424	: data2 <= weights[3425];
				12'd3425	: data2 <= weights[3426];
				12'd3426	: data2 <= weights[3427];
				12'd3427	: data2 <= weights[3428];
				12'd3428	: data2 <= weights[3429];
				12'd3429	: data2 <= weights[3430];
				12'd3430	: data2 <= weights[3431];
				12'd3431	: data2 <= weights[3432];
				12'd3432	: data2 <= weights[3433];
				12'd3433	: data2 <= weights[3434];
				12'd3434	: data2 <= weights[3435];
				12'd3435	: data2 <= weights[3436];
				12'd3436	: data2 <= weights[3437];
				12'd3437	: data2 <= weights[3438];
				12'd3438	: data2 <= weights[3439];
				12'd3439	: data2 <= weights[3440];
				12'd3440	: data2 <= weights[3441];
				12'd3441	: data2 <= weights[3442];
				12'd3442	: data2 <= weights[3443];
				12'd3443	: data2 <= weights[3444];
				12'd3444	: data2 <= weights[3445];
				12'd3445	: data2 <= weights[3446];
				12'd3446	: data2 <= weights[3447];
				12'd3447	: data2 <= weights[3448];
				12'd3448	: data2 <= weights[3449];
				12'd3449	: data2 <= weights[3450];
				12'd3450	: data2 <= weights[3451];
				12'd3451	: data2 <= weights[3452];
				12'd3452	: data2 <= weights[3453];
				12'd3453	: data2 <= weights[3454];
				12'd3454	: data2 <= weights[3455];
				12'd3455	: data2 <= weights[3456];
				12'd3456	: data2 <= weights[3457];
				12'd3457	: data2 <= weights[3458];
				12'd3458	: data2 <= weights[3459];
				12'd3459	: data2 <= weights[3460];
				12'd3460	: data2 <= weights[3461];
				12'd3461	: data2 <= weights[3462];
				12'd3462	: data2 <= weights[3463];
				12'd3463	: data2 <= weights[3464];
				12'd3464	: data2 <= weights[3465];
				12'd3465	: data2 <= weights[3466];
				12'd3466	: data2 <= weights[3467];
				12'd3467	: data2 <= weights[3468];
				12'd3468	: data2 <= weights[3469];
				12'd3469	: data2 <= weights[3470];
				12'd3470	: data2 <= weights[3471];
				12'd3471	: data2 <= weights[3472];
				12'd3472	: data2 <= weights[3473];
				12'd3473	: data2 <= weights[3474];
				12'd3474	: data2 <= weights[3475];
				12'd3475	: data2 <= weights[3476];
				12'd3476	: data2 <= weights[3477];
				12'd3477	: data2 <= weights[3478];
				12'd3478	: data2 <= weights[3479];
				12'd3479	: data2 <= weights[3480];
				12'd3480	: data2 <= weights[3481];
				12'd3481	: data2 <= weights[3482];
				12'd3482	: data2 <= weights[3483];
				12'd3483	: data2 <= weights[3484];
				12'd3484	: data2 <= weights[3485];
				12'd3485	: data2 <= weights[3486];
				12'd3486	: data2 <= weights[3487];
				12'd3487	: data2 <= weights[3488];
				12'd3488	: data2 <= weights[3489];
				12'd3489	: data2 <= weights[3490];
				12'd3490	: data2 <= weights[3491];
				12'd3491	: data2 <= weights[3492];
				12'd3492	: data2 <= weights[3493];
				12'd3493	: data2 <= weights[3494];
				12'd3494	: data2 <= weights[3495];
				12'd3495	: data2 <= weights[3496];
				12'd3496	: data2 <= weights[3497];
				12'd3497	: data2 <= weights[3498];
				12'd3498	: data2 <= weights[3499];
				12'd3499	: data2 <= weights[3500];
				12'd3500	: data2 <= weights[3501];
				12'd3501	: data2 <= weights[3502];
				12'd3502	: data2 <= weights[3503];
				12'd3503	: data2 <= weights[3504];
				12'd3504	: data2 <= weights[3505];
				12'd3505	: data2 <= weights[3506];
				12'd3506	: data2 <= weights[3507];
				12'd3507	: data2 <= weights[3508];
				12'd3508	: data2 <= weights[3509];
				12'd3509	: data2 <= weights[3510];
				12'd3510	: data2 <= weights[3511];
				12'd3511	: data2 <= weights[3512];
				12'd3512	: data2 <= weights[3513];
				12'd3513	: data2 <= weights[3514];
				12'd3514	: data2 <= weights[3515];
				12'd3515	: data2 <= weights[3516];
				12'd3516	: data2 <= weights[3517];
				12'd3517	: data2 <= weights[3518];
				12'd3518	: data2 <= weights[3519];
				12'd3519	: data2 <= weights[3520];
				12'd3520	: data2 <= weights[3521];
				12'd3521	: data2 <= weights[3522];
				12'd3522	: data2 <= weights[3523];
				12'd3523	: data2 <= weights[3524];
				12'd3524	: data2 <= weights[3525];
				12'd3525	: data2 <= weights[3526];
				12'd3526	: data2 <= weights[3527];
				12'd3527	: data2 <= weights[3528];
				12'd3528	: data2 <= weights[3529];
				12'd3529	: data2 <= weights[3530];
				12'd3530	: data2 <= weights[3531];
				12'd3531	: data2 <= weights[3532];
				12'd3532	: data2 <= weights[3533];
				12'd3533	: data2 <= weights[3534];
				12'd3534	: data2 <= weights[3535];
				12'd3535	: data2 <= weights[3536];
				12'd3536	: data2 <= weights[3537];
				12'd3537	: data2 <= weights[3538];
				12'd3538	: data2 <= weights[3539];
				12'd3539	: data2 <= weights[3540];
				12'd3540	: data2 <= weights[3541];
				12'd3541	: data2 <= weights[3542];
				12'd3542	: data2 <= weights[3543];
				12'd3543	: data2 <= weights[3544];
				12'd3544	: data2 <= weights[3545];
				12'd3545	: data2 <= weights[3546];
				12'd3546	: data2 <= weights[3547];
				12'd3547	: data2 <= weights[3548];
				12'd3548	: data2 <= weights[3549];
				12'd3549	: data2 <= weights[3550];
				12'd3550	: data2 <= weights[3551];
				12'd3551	: data2 <= weights[3552];
				12'd3552	: data2 <= weights[3553];
				12'd3553	: data2 <= weights[3554];
				12'd3554	: data2 <= weights[3555];
				12'd3555	: data2 <= weights[3556];
				12'd3556	: data2 <= weights[3557];
				12'd3557	: data2 <= weights[3558];
				12'd3558	: data2 <= weights[3559];
				12'd3559	: data2 <= weights[3560];
				12'd3560	: data2 <= weights[3561];
				12'd3561	: data2 <= weights[3562];
				12'd3562	: data2 <= weights[3563];
				12'd3563	: data2 <= weights[3564];
				12'd3564	: data2 <= weights[3565];
				12'd3565	: data2 <= weights[3566];
				12'd3566	: data2 <= weights[3567];
				12'd3567	: data2 <= weights[3568];
				12'd3568	: data2 <= weights[3569];
				12'd3569	: data2 <= weights[3570];
				12'd3570	: data2 <= weights[3571];
				12'd3571	: data2 <= weights[3572];
				12'd3572	: data2 <= weights[3573];
				12'd3573	: data2 <= weights[3574];
				12'd3574	: data2 <= weights[3575];
				12'd3575	: data2 <= weights[3576];
				12'd3576	: data2 <= weights[3577];
				12'd3577	: data2 <= weights[3578];
				12'd3578	: data2 <= weights[3579];
				12'd3579	: data2 <= weights[3580];
				12'd3580	: data2 <= weights[3581];
				12'd3581	: data2 <= weights[3582];
				12'd3582	: data2 <= weights[3583];
				12'd3583	: data2 <= weights[3584];
				12'd3584	: data2 <= weights[3585];
				12'd3585	: data2 <= weights[3586];
				12'd3586	: data2 <= weights[3587];
				12'd3587	: data2 <= weights[3588];
				12'd3588	: data2 <= weights[3589];
				12'd3589	: data2 <= weights[3590];
				12'd3590	: data2 <= weights[3591];
				12'd3591	: data2 <= weights[3592];
				12'd3592	: data2 <= weights[3593];
				12'd3593	: data2 <= weights[3594];
				12'd3594	: data2 <= weights[3595];
				12'd3595	: data2 <= weights[3596];
				12'd3596	: data2 <= weights[3597];
				12'd3597	: data2 <= weights[3598];
				12'd3598	: data2 <= weights[3599];
				12'd3599	: data2 <= weights[3600];
				12'd3600	: data2 <= weights[3601];
				12'd3601	: data2 <= weights[3602];
				12'd3602	: data2 <= weights[3603];
				12'd3603	: data2 <= weights[3604];
				12'd3604	: data2 <= weights[3605];
				12'd3605	: data2 <= weights[3606];
				12'd3606	: data2 <= weights[3607];
				12'd3607	: data2 <= weights[3608];
				12'd3608	: data2 <= weights[3609];
				12'd3609	: data2 <= weights[3610];
				12'd3610	: data2 <= weights[3611];
				12'd3611	: data2 <= weights[3612];
				12'd3612	: data2 <= weights[3613];
				12'd3613	: data2 <= weights[3614];
				12'd3614	: data2 <= weights[3615];
				12'd3615	: data2 <= weights[3616];
				12'd3616	: data2 <= weights[3617];
				12'd3617	: data2 <= weights[3618];
				12'd3618	: data2 <= weights[3619];
				12'd3619	: data2 <= weights[3620];
				12'd3620	: data2 <= weights[3621];
				12'd3621	: data2 <= weights[3622];
				12'd3622	: data2 <= weights[3623];
				12'd3623	: data2 <= weights[3624];
				12'd3624	: data2 <= weights[3625];
				12'd3625	: data2 <= weights[3626];
				12'd3626	: data2 <= weights[3627];
				12'd3627	: data2 <= weights[3628];
				12'd3628	: data2 <= weights[3629];
				12'd3629	: data2 <= weights[3630];
				12'd3630	: data2 <= weights[3631];
				12'd3631	: data2 <= weights[3632];
				12'd3632	: data2 <= weights[3633];
				12'd3633	: data2 <= weights[3634];
				12'd3634	: data2 <= weights[3635];
				12'd3635	: data2 <= weights[3636];
				12'd3636	: data2 <= weights[3637];
				12'd3637	: data2 <= weights[3638];
				12'd3638	: data2 <= weights[3639];
				12'd3639	: data2 <= weights[3640];
				12'd3640	: data2 <= weights[3641];
				12'd3641	: data2 <= weights[3642];
				12'd3642	: data2 <= weights[3643];
				12'd3643	: data2 <= weights[3644];
				12'd3644	: data2 <= weights[3645];
				12'd3645	: data2 <= weights[3646];
				12'd3646	: data2 <= weights[3647];
				12'd3647	: data2 <= weights[3648];
				12'd3648	: data2 <= weights[3649];
				12'd3649	: data2 <= weights[3650];
				12'd3650	: data2 <= weights[3651];
				12'd3651	: data2 <= weights[3652];
				12'd3652	: data2 <= weights[3653];
				12'd3653	: data2 <= weights[3654];
				12'd3654	: data2 <= weights[3655];
				12'd3655	: data2 <= weights[3656];
				12'd3656	: data2 <= weights[3657];
				12'd3657	: data2 <= weights[3658];
				12'd3658	: data2 <= weights[3659];
				12'd3659	: data2 <= weights[3660];
				12'd3660	: data2 <= weights[3661];
				12'd3661	: data2 <= weights[3662];
				12'd3662	: data2 <= weights[3663];
				12'd3663	: data2 <= weights[3664];
				12'd3664	: data2 <= weights[3665];
				12'd3665	: data2 <= weights[3666];
				12'd3666	: data2 <= weights[3667];
				12'd3667	: data2 <= weights[3668];
				12'd3668	: data2 <= weights[3669];
				12'd3669	: data2 <= weights[3670];
				12'd3670	: data2 <= weights[3671];
				12'd3671	: data2 <= weights[3672];
				12'd3672	: data2 <= weights[3673];
				12'd3673	: data2 <= weights[3674];
				12'd3674	: data2 <= weights[3675];
				12'd3675	: data2 <= weights[3676];
				12'd3676	: data2 <= weights[3677];
				12'd3677	: data2 <= weights[3678];
				12'd3678	: data2 <= weights[3679];
				12'd3679	: data2 <= weights[3680];
				12'd3680	: data2 <= weights[3681];
				12'd3681	: data2 <= weights[3682];
				12'd3682	: data2 <= weights[3683];
				12'd3683	: data2 <= weights[3684];
				12'd3684	: data2 <= weights[3685];
				12'd3685	: data2 <= weights[3686];
				12'd3686	: data2 <= weights[3687];
				12'd3687	: data2 <= weights[3688];
				12'd3688	: data2 <= weights[3689];
				12'd3689	: data2 <= weights[3690];
				12'd3690	: data2 <= weights[3691];
				12'd3691	: data2 <= weights[3692];
				12'd3692	: data2 <= weights[3693];
				12'd3693	: data2 <= weights[3694];
				12'd3694	: data2 <= weights[3695];
				12'd3695	: data2 <= weights[3696];
				12'd3696	: data2 <= weights[3697];
				12'd3697	: data2 <= weights[3698];
				12'd3698	: data2 <= weights[3699];
				12'd3699	: data2 <= weights[3700];
				12'd3700	: data2 <= weights[3701];
				12'd3701	: data2 <= weights[3702];
				12'd3702	: data2 <= weights[3703];
				12'd3703	: data2 <= weights[3704];
				12'd3704	: data2 <= weights[3705];
				12'd3705	: data2 <= weights[3706];
				12'd3706	: data2 <= weights[3707];
				12'd3707	: data2 <= weights[3708];
				12'd3708	: data2 <= weights[3709];
				12'd3709	: data2 <= weights[3710];
				12'd3710	: data2 <= weights[3711];
				12'd3711	: data2 <= weights[3712];
				12'd3712	: data2 <= weights[3713];
				12'd3713	: data2 <= weights[3714];
				12'd3714	: data2 <= weights[3715];
				12'd3715	: data2 <= weights[3716];
				12'd3716	: data2 <= weights[3717];
				12'd3717	: data2 <= weights[3718];
				12'd3718	: data2 <= weights[3719];
				12'd3719	: data2 <= weights[3720];
				12'd3720	: data2 <= weights[3721];
				12'd3721	: data2 <= weights[3722];
				12'd3722	: data2 <= weights[3723];
				12'd3723	: data2 <= weights[3724];
				12'd3724	: data2 <= weights[3725];
				12'd3725	: data2 <= weights[3726];
				12'd3726	: data2 <= weights[3727];
				12'd3727	: data2 <= weights[3728];
				12'd3728	: data2 <= weights[3729];
				12'd3729	: data2 <= weights[3730];
				12'd3730	: data2 <= weights[3731];
				12'd3731	: data2 <= weights[3732];
				12'd3732	: data2 <= weights[3733];
				12'd3733	: data2 <= weights[3734];
				12'd3734	: data2 <= weights[3735];
				12'd3735	: data2 <= weights[3736];
				12'd3736	: data2 <= weights[3737];
				12'd3737	: data2 <= weights[3738];
				12'd3738	: data2 <= weights[3739];
				12'd3739	: data2 <= weights[3740];
				12'd3740	: data2 <= weights[3741];
				12'd3741	: data2 <= weights[3742];
				12'd3742	: data2 <= weights[3743];
				12'd3743	: data2 <= weights[3744];
				12'd3744	: data2 <= weights[3745];
				12'd3745	: data2 <= weights[3746];
				12'd3746	: data2 <= weights[3747];
				12'd3747	: data2 <= weights[3748];
				12'd3748	: data2 <= weights[3749];
				12'd3749	: data2 <= weights[3750];
				12'd3750	: data2 <= weights[3751];
				12'd3751	: data2 <= weights[3752];
				12'd3752	: data2 <= weights[3753];
				12'd3753	: data2 <= weights[3754];
				12'd3754	: data2 <= weights[3755];
				12'd3755	: data2 <= weights[3756];
				12'd3756	: data2 <= weights[3757];
				12'd3757	: data2 <= weights[3758];
				12'd3758	: data2 <= weights[3759];
				12'd3759	: data2 <= weights[3760];
				12'd3760	: data2 <= weights[3761];
				12'd3761	: data2 <= weights[3762];
				12'd3762	: data2 <= weights[3763];
				12'd3763	: data2 <= weights[3764];
				12'd3764	: data2 <= weights[3765];
				12'd3765	: data2 <= weights[3766];
				12'd3766	: data2 <= weights[3767];
				12'd3767	: data2 <= weights[3768];
				12'd3768	: data2 <= weights[3769];
				12'd3769	: data2 <= weights[3770];
				12'd3770	: data2 <= weights[3771];
				12'd3771	: data2 <= weights[3772];
				12'd3772	: data2 <= weights[3773];
				12'd3773	: data2 <= weights[3774];
				12'd3774	: data2 <= weights[3775];
				12'd3775	: data2 <= weights[3776];
				12'd3776	: data2 <= weights[3777];
				12'd3777	: data2 <= weights[3778];
				12'd3778	: data2 <= weights[3779];
				12'd3779	: data2 <= weights[3780];
				12'd3780	: data2 <= weights[3781];
				12'd3781	: data2 <= weights[3782];
				12'd3782	: data2 <= weights[3783];
				12'd3783	: data2 <= weights[3784];
				12'd3784	: data2 <= weights[3785];
				12'd3785	: data2 <= weights[3786];
				12'd3786	: data2 <= weights[3787];
				12'd3787	: data2 <= weights[3788];
				12'd3788	: data2 <= weights[3789];
				12'd3789	: data2 <= weights[3790];
				12'd3790	: data2 <= weights[3791];
				12'd3791	: data2 <= weights[3792];
				12'd3792	: data2 <= weights[3793];
				12'd3793	: data2 <= weights[3794];
				12'd3794	: data2 <= weights[3795];
				12'd3795	: data2 <= weights[3796];
				12'd3796	: data2 <= weights[3797];
				12'd3797	: data2 <= weights[3798];
				12'd3798	: data2 <= weights[3799];
				12'd3799	: data2 <= weights[3800];
				12'd3800	: data2 <= weights[3801];
				12'd3801	: data2 <= weights[3802];
				12'd3802	: data2 <= weights[3803];
				12'd3803	: data2 <= weights[3804];
				12'd3804	: data2 <= weights[3805];
				12'd3805	: data2 <= weights[3806];
				12'd3806	: data2 <= weights[3807];
				12'd3807	: data2 <= weights[3808];
				12'd3808	: data2 <= weights[3809];
				12'd3809	: data2 <= weights[3810];
				12'd3810	: data2 <= weights[3811];
				12'd3811	: data2 <= weights[3812];
				12'd3812	: data2 <= weights[3813];
				12'd3813	: data2 <= weights[3814];
				12'd3814	: data2 <= weights[3815];
				12'd3815	: data2 <= weights[3816];
				12'd3816	: data2 <= weights[3817];
				12'd3817	: data2 <= weights[3818];
				12'd3818	: data2 <= weights[3819];
				12'd3819	: data2 <= weights[3820];
				12'd3820	: data2 <= weights[3821];
				12'd3821	: data2 <= weights[3822];
				12'd3822	: data2 <= weights[3823];
				12'd3823	: data2 <= weights[3824];
				12'd3824	: data2 <= weights[3825];
				12'd3825	: data2 <= weights[3826];
				12'd3826	: data2 <= weights[3827];
				12'd3827	: data2 <= weights[3828];
				12'd3828	: data2 <= weights[3829];
				12'd3829	: data2 <= weights[3830];
				12'd3830	: data2 <= weights[3831];
				12'd3831	: data2 <= weights[3832];
				12'd3832	: data2 <= weights[3833];
				12'd3833	: data2 <= weights[3834];
				12'd3834	: data2 <= weights[3835];
				12'd3835	: data2 <= weights[3836];
				12'd3836	: data2 <= weights[3837];
				12'd3837	: data2 <= weights[3838];
				12'd3838	: data2 <= weights[3839];
				12'd3839	: data2 <= weights[3840];
				12'd3840	: data2 <= weights[3841];
				12'd3841	: data2 <= weights[3842];
				12'd3842	: data2 <= weights[3843];
				12'd3843	: data2 <= weights[3844];
				12'd3844	: data2 <= weights[3845];
				12'd3845	: data2 <= weights[3846];
				12'd3846	: data2 <= weights[3847];
				12'd3847	: data2 <= weights[3848];
				12'd3848	: data2 <= weights[3849];
				12'd3849	: data2 <= weights[3850];
				12'd3850	: data2 <= weights[3851];
				12'd3851	: data2 <= weights[3852];
				12'd3852	: data2 <= weights[3853];
				12'd3853	: data2 <= weights[3854];
				12'd3854	: data2 <= weights[3855];
				12'd3855	: data2 <= weights[3856];
				12'd3856	: data2 <= weights[3857];
				12'd3857	: data2 <= weights[3858];
				12'd3858	: data2 <= weights[3859];
				12'd3859	: data2 <= weights[3860];
				12'd3860	: data2 <= weights[3861];
				12'd3861	: data2 <= weights[3862];
				12'd3862	: data2 <= weights[3863];
				12'd3863	: data2 <= weights[3864];
				12'd3864	: data2 <= weights[3865];
				12'd3865	: data2 <= weights[3866];
				12'd3866	: data2 <= weights[3867];
				12'd3867	: data2 <= weights[3868];
				12'd3868	: data2 <= weights[3869];
				12'd3869	: data2 <= weights[3870];
				12'd3870	: data2 <= weights[3871];
				12'd3871	: data2 <= weights[3872];
				12'd3872	: data2 <= weights[3873];
				12'd3873	: data2 <= weights[3874];
				12'd3874	: data2 <= weights[3875];
				12'd3875	: data2 <= weights[3876];
				12'd3876	: data2 <= weights[3877];
				12'd3877	: data2 <= weights[3878];
				12'd3878	: data2 <= weights[3879];
				12'd3879	: data2 <= weights[3880];
				12'd3880	: data2 <= weights[3881];
				12'd3881	: data2 <= weights[3882];
				12'd3882	: data2 <= weights[3883];
				12'd3883	: data2 <= weights[3884];
				12'd3884	: data2 <= weights[3885];
				12'd3885	: data2 <= weights[3886];
				12'd3886	: data2 <= weights[3887];
				12'd3887	: data2 <= weights[3888];
				12'd3888	: data2 <= weights[3889];
				12'd3889	: data2 <= weights[3890];
				12'd3890	: data2 <= weights[3891];
				12'd3891	: data2 <= weights[3892];
				12'd3892	: data2 <= weights[3893];
				12'd3893	: data2 <= weights[3894];
				12'd3894	: data2 <= weights[3895];
				12'd3895	: data2 <= weights[3896];
				12'd3896	: data2 <= weights[3897];
				12'd3897	: data2 <= weights[3898];
				12'd3898	: data2 <= weights[3899];
				12'd3899	: data2 <= weights[3900];
				12'd3900	: data2 <= weights[3901];
				12'd3901	: data2 <= weights[3902];
				12'd3902	: data2 <= weights[3903];
				12'd3903	: data2 <= weights[3904];
				12'd3904	: data2 <= weights[3905];
				12'd3905	: data2 <= weights[3906];
				12'd3906	: data2 <= weights[3907];
				12'd3907	: data2 <= weights[3908];
				12'd3908	: data2 <= weights[3909];
				12'd3909	: data2 <= weights[3910];
				12'd3910	: data2 <= weights[3911];
				12'd3911	: data2 <= weights[3912];
				12'd3912	: data2 <= weights[3913];
				12'd3913	: data2 <= weights[3914];
				12'd3914	: data2 <= weights[3915];
				12'd3915	: data2 <= weights[3916];
				12'd3916	: data2 <= weights[3917];
				12'd3917	: data2 <= weights[3918];
				12'd3918	: data2 <= weights[3919];
				12'd3919	: data2 <= weights[3920];
				12'd3920	: data2 <= weights[3921];
				12'd3921	: data2 <= weights[3922];
				12'd3922	: data2 <= weights[3923];
				12'd3923	: data2 <= weights[3924];
				12'd3924	: data2 <= weights[3925];
				12'd3925	: data2 <= weights[3926];
				12'd3926	: data2 <= weights[3927];
				12'd3927	: data2 <= weights[3928];
				12'd3928	: data2 <= weights[3929];
				12'd3929	: data2 <= weights[3930];
				12'd3930	: data2 <= weights[3931];
				12'd3931	: data2 <= weights[3932];
				12'd3932	: data2 <= weights[3933];
				12'd3933	: data2 <= weights[3934];
				12'd3934	: data2 <= weights[3935];
				12'd3935	: data2 <= weights[3936];
				12'd3936	: data2 <= weights[3937];
				12'd3937	: data2 <= weights[3938];
				12'd3938	: data2 <= weights[3939];
				12'd3939	: data2 <= weights[3940];
				12'd3940	: data2 <= weights[3941];
				12'd3941	: data2 <= weights[3942];
				12'd3942	: data2 <= weights[3943];
				12'd3943	: data2 <= weights[3944];
				12'd3944	: data2 <= weights[3945];
				12'd3945	: data2 <= weights[3946];
				12'd3946	: data2 <= weights[3947];
				12'd3947	: data2 <= weights[3948];
				12'd3948	: data2 <= weights[3949];
				12'd3949	: data2 <= weights[3950];
				12'd3950	: data2 <= weights[3951];
				12'd3951	: data2 <= weights[3952];
				12'd3952	: data2 <= weights[3953];
				12'd3953	: data2 <= weights[3954];
				12'd3954	: data2 <= weights[3955];
				12'd3955	: data2 <= weights[3956];
				12'd3956	: data2 <= weights[3957];
				12'd3957	: data2 <= weights[3958];
				12'd3958	: data2 <= weights[3959];
				12'd3959	: data2 <= weights[3960];
				12'd3960	: data2 <= weights[3961];
				12'd3961	: data2 <= weights[3962];
				12'd3962	: data2 <= weights[3963];
				12'd3963	: data2 <= weights[3964];
				12'd3964	: data2 <= weights[3965];
				12'd3965	: data2 <= weights[3966];
				12'd3966	: data2 <= weights[3967];
				12'd3967	: data2 <= weights[3968];
				12'd3968	: data2 <= weights[3969];
				12'd3969	: data2 <= weights[3970];
				12'd3970	: data2 <= weights[3971];
				12'd3971	: data2 <= weights[3972];
				12'd3972	: data2 <= weights[3973];
				12'd3973	: data2 <= weights[3974];
				12'd3974	: data2 <= weights[3975];
				12'd3975	: data2 <= weights[3976];
				12'd3976	: data2 <= weights[3977];
				12'd3977	: data2 <= weights[3978];
				12'd3978	: data2 <= weights[3979];
				12'd3979	: data2 <= weights[3980];
				12'd3980	: data2 <= weights[3981];
				12'd3981	: data2 <= weights[3982];
				12'd3982	: data2 <= weights[3983];
				12'd3983	: data2 <= weights[3984];
				12'd3984	: data2 <= weights[3985];
				12'd3985	: data2 <= weights[3986];
				12'd3986	: data2 <= weights[3987];
				12'd3987	: data2 <= weights[3988];
				12'd3988	: data2 <= weights[3989];
				12'd3989	: data2 <= weights[3990];
				12'd3990	: data2 <= weights[3991];
				12'd3991	: data2 <= weights[3992];
				12'd3992	: data2 <= weights[3993];
				12'd3993	: data2 <= weights[3994];
				12'd3994	: data2 <= weights[3995];
				12'd3995	: data2 <= weights[3996];
				12'd3996	: data2 <= weights[3997];
				12'd3997	: data2 <= weights[3998];
				12'd3998	: data2 <= weights[3999];
				12'd3999	: data2 <= weights[4000];
				12'd4000	: data2 <= weights[4001];
				12'd4001	: data2 <= weights[4002];
				12'd4002	: data2 <= weights[4003];
				12'd4003	: data2 <= weights[4004];
				12'd4004	: data2 <= weights[4005];
				12'd4005	: data2 <= weights[4006];
				12'd4006	: data2 <= weights[4007];
				12'd4007	: data2 <= weights[4008];
				12'd4008	: data2 <= weights[4009];
				12'd4009	: data2 <= weights[4010];
				12'd4010	: data2 <= weights[4011];
				12'd4011	: data2 <= weights[4012];
				12'd4012	: data2 <= weights[4013];
				12'd4013	: data2 <= weights[4014];
				12'd4014	: data2 <= weights[4015];
				12'd4015	: data2 <= weights[4016];
				12'd4016	: data2 <= weights[4017];
				12'd4017	: data2 <= weights[4018];
				12'd4018	: data2 <= weights[4019];
				12'd4019	: data2 <= weights[4020];
				12'd4020	: data2 <= weights[4021];
				12'd4021	: data2 <= weights[4022];
				12'd4022	: data2 <= weights[4023];
				12'd4023	: data2 <= weights[4024];
				12'd4024	: data2 <= weights[4025];
				12'd4025	: data2 <= weights[4026];
				12'd4026	: data2 <= weights[4027];
				12'd4027	: data2 <= weights[4028];
				12'd4028	: data2 <= weights[4029];
				12'd4029	: data2 <= weights[4030];
				12'd4030	: data2 <= weights[4031];
				12'd4031	: data2 <= weights[4032];
				12'd4032	: data2 <= weights[4033];
				12'd4033	: data2 <= weights[4034];
				12'd4034	: data2 <= weights[4035];
				12'd4035	: data2 <= weights[4036];
				12'd4036	: data2 <= weights[4037];
				12'd4037	: data2 <= weights[4038];
				12'd4038	: data2 <= weights[4039];
				12'd4039	: data2 <= weights[4040];
				12'd4040	: data2 <= weights[4041];
				12'd4041	: data2 <= weights[4042];
				12'd4042	: data2 <= weights[4043];
				12'd4043	: data2 <= weights[4044];
				12'd4044	: data2 <= weights[4045];
				12'd4045	: data2 <= weights[4046];
				12'd4046	: data2 <= weights[4047];
				12'd4047	: data2 <= weights[4048];
				12'd4048	: data2 <= weights[4049];
				12'd4049	: data2 <= weights[4050];
				default		: data2 <= 16'd0;
			endcase
		end else begin
			data2 <= data2;
		end
	end

endmodule