module ROM(
	input wire clk,
	input wire enable,
	input wire [11:0] address,
	output reg [15:0] data1,
	output reg [15:0] data2
	);

	reg [15:0] weights [4050:0];

	initial begin
		weights[0] <= 171;
		weights[1] <= 189;
		weights[2] <= 109;
		weights[3] <= 186;
		weights[4] <= 71;
		weights[5] <= 46;
		weights[6] <= 170;
		weights[7] <= 91;
		weights[8] <= 251;
		weights[9] <= 56;
		weights[10] <= 3;
		weights[11] <= 145;
		weights[12] <= 100;
		weights[13] <= 38;
		weights[14] <= 74;
		weights[15] <= 137;
		weights[16] <= 80;
		weights[17] <= 19;
		weights[18] <= 185;
		weights[19] <= 177;
		weights[20] <= 178;
		weights[21] <= 222;
		weights[22] <= 201;
		weights[23] <= 107;
		weights[24] <= 202;
		weights[25] <= 171;
		weights[26] <= 216;
		weights[27] <= 94;
		weights[28] <= 95;
		weights[29] <= 190;
		weights[30] <= 9;
		weights[31] <= 230;
		weights[32] <= 80;
		weights[33] <= 26;
		weights[34] <= 225;
		weights[35] <= 19;
		weights[36] <= 29;
		weights[37] <= 61;
		weights[38] <= 93;
		weights[39] <= 253;
		weights[40] <= 83;
		weights[41] <= 201;
		weights[42] <= 226;
		weights[43] <= 113;
		weights[44] <= 145;
		weights[45] <= 144;
		weights[46] <= 84;
		weights[47] <= 185;
		weights[48] <= 179;
		weights[49] <= 141;
		weights[50] <= 226;
		weights[51] <= 142;
		weights[52] <= 169;
		weights[53] <= 17;
		weights[54] <= 153;
		weights[55] <= 249;
		weights[56] <= 82;
		weights[57] <= 95;
		weights[58] <= 163;
		weights[59] <= 146;
		weights[60] <= 94;
		weights[61] <= 22;
		weights[62] <= 11;
		weights[63] <= 205;
		weights[64] <= 186;
		weights[65] <= 209;
		weights[66] <= 243;
		weights[67] <= 127;
		weights[68] <= 59;
		weights[69] <= 66;
		weights[70] <= 223;
		weights[71] <= 79;
		weights[72] <= 247;
		weights[73] <= 34;
		weights[74] <= 25;
		weights[75] <= 91;
		weights[76] <= 81;
		weights[77] <= 253;
		weights[78] <= 6;
		weights[79] <= 168;
		weights[80] <= 192;
		weights[81] <= 26;
		weights[82] <= 250;
		weights[83] <= 82;
		weights[84] <= 247;
		weights[85] <= 39;
		weights[86] <= 212;
		weights[87] <= 127;
		weights[88] <= 144;
		weights[89] <= 178;
		weights[90] <= 165;
		weights[91] <= 89;
		weights[92] <= 38;
		weights[93] <= 221;
		weights[94] <= 253;
		weights[95] <= 210;
		weights[96] <= 248;
		weights[97] <= 246;
		weights[98] <= 162;
		weights[99] <= 87;
		weights[100] <= 85;
		weights[101] <= 19;
		weights[102] <= 164;
		weights[103] <= 213;
		weights[104] <= 80;
		weights[105] <= 236;
		weights[106] <= 93;
		weights[107] <= 179;
		weights[108] <= 197;
		weights[109] <= 45;
		weights[110] <= 141;
		weights[111] <= 88;
		weights[112] <= 183;
		weights[113] <= 114;
		weights[114] <= 203;
		weights[115] <= 121;
		weights[116] <= 31;
		weights[117] <= 180;
		weights[118] <= 146;
		weights[119] <= 247;
		weights[120] <= 246;
		weights[121] <= 102;
		weights[122] <= 32;
		weights[123] <= 225;
		weights[124] <= 37;
		weights[125] <= 222;
		weights[126] <= 216;
		weights[127] <= 195;
		weights[128] <= 182;
		weights[129] <= 203;
		weights[130] <= 43;
		weights[131] <= 72;
		weights[132] <= 229;
		weights[133] <= 172;
		weights[134] <= 202;
		weights[135] <= 56;
		weights[136] <= 72;
		weights[137] <= 131;
		weights[138] <= 16;
		weights[139] <= 51;
		weights[140] <= 99;
		weights[141] <= 54;
		weights[142] <= 196;
		weights[143] <= 163;
		weights[144] <= 195;
		weights[145] <= 112;
		weights[146] <= 95;
		weights[147] <= 63;
		weights[148] <= 228;
		weights[149] <= 16;
		weights[150] <= 239;
		weights[151] <= 107;
		weights[152] <= 32;
		weights[153] <= 117;
		weights[154] <= 154;
		weights[155] <= 48;
		weights[156] <= 2;
		weights[157] <= 11;
		weights[158] <= 109;
		weights[159] <= 95;
		weights[160] <= 117;
		weights[161] <= 183;
		weights[162] <= 111;
		weights[163] <= 5;
		weights[164] <= 212;
		weights[165] <= 32;
		weights[166] <= 201;
		weights[167] <= 63;
		weights[168] <= 165;
		weights[169] <= 43;
		weights[170] <= 233;
		weights[171] <= 238;
		weights[172] <= 25;
		weights[173] <= 36;
		weights[174] <= 250;
		weights[175] <= 200;
		weights[176] <= 218;
		weights[177] <= 145;
		weights[178] <= 135;
		weights[179] <= 207;
		weights[180] <= 201;
		weights[181] <= 107;
		weights[182] <= 204;
		weights[183] <= 12;
		weights[184] <= 219;
		weights[185] <= 238;
		weights[186] <= 253;
		weights[187] <= 252;
		weights[188] <= 225;
		weights[189] <= 247;
		weights[190] <= 196;
		weights[191] <= 197;
		weights[192] <= 234;
		weights[193] <= 189;
		weights[194] <= 166;
		weights[195] <= 27;
		weights[196] <= 10;
		weights[197] <= 91;
		weights[198] <= 163;
		weights[199] <= 190;
		weights[200] <= 63;
		weights[201] <= 228;
		weights[202] <= 64;
		weights[203] <= 172;
		weights[204] <= 191;
		weights[205] <= 198;
		weights[206] <= 155;
		weights[207] <= 152;
		weights[208] <= 165;
		weights[209] <= 233;
		weights[210] <= 250;
		weights[211] <= 250;
		weights[212] <= 16;
		weights[213] <= 247;
		weights[214] <= 57;
		weights[215] <= 46;
		weights[216] <= 241;
		weights[217] <= 230;
		weights[218] <= 244;
		weights[219] <= 182;
		weights[220] <= 58;
		weights[221] <= 253;
		weights[222] <= 115;
		weights[223] <= 166;
		weights[224] <= 81;
		weights[225] <= 161;
		weights[226] <= 223;
		weights[227] <= 220;
		weights[228] <= 25;
		weights[229] <= 118;
		weights[230] <= 162;
		weights[231] <= 42;
		weights[232] <= 237;
		weights[233] <= 218;
		weights[234] <= 198;
		weights[235] <= 200;
		weights[236] <= 80;
		weights[237] <= 150;
		weights[238] <= 156;
		weights[239] <= 80;
		weights[240] <= 102;
		weights[241] <= 32;
		weights[242] <= 22;
		weights[243] <= 21;
		weights[244] <= 222;
		weights[245] <= 217;
		weights[246] <= 193;
		weights[247] <= 244;
		weights[248] <= 88;
		weights[249] <= 46;
		weights[250] <= 50;
		weights[251] <= 211;
		weights[252] <= 218;
		weights[253] <= 228;
		weights[254] <= 250;
		weights[255] <= 137;
		weights[256] <= 66;
		weights[257] <= 194;
		weights[258] <= 203;
		weights[259] <= 120;
		weights[260] <= 79;
		weights[261] <= 118;
		weights[262] <= 60;
		weights[263] <= 220;
		weights[264] <= 32;
		weights[265] <= 55;
		weights[266] <= 143;
		weights[267] <= 15;
		weights[268] <= 255;
		weights[269] <= 128;
		weights[270] <= 123;
		weights[271] <= 238;
		weights[272] <= 55;
		weights[273] <= 14;
		weights[274] <= 240;
		weights[275] <= 136;
		weights[276] <= 77;
		weights[277] <= 130;
		weights[278] <= 74;
		weights[279] <= 9;
		weights[280] <= 201;
		weights[281] <= 156;
		weights[282] <= 94;
		weights[283] <= 124;
		weights[284] <= 36;
		weights[285] <= 27;
		weights[286] <= 51;
		weights[287] <= 196;
		weights[288] <= 86;
		weights[289] <= 23;
		weights[290] <= 92;
		weights[291] <= 17;
		weights[292] <= 133;
		weights[293] <= 139;
		weights[294] <= 229;
		weights[295] <= 13;
		weights[296] <= 209;
		weights[297] <= 75;
		weights[298] <= 134;
		weights[299] <= 210;
		weights[300] <= 156;
		weights[301] <= 142;
		weights[302] <= 206;
		weights[303] <= 122;
		weights[304] <= 155;
		weights[305] <= 122;
		weights[306] <= 29;
		weights[307] <= 77;
		weights[308] <= 80;
		weights[309] <= 74;
		weights[310] <= 69;
		weights[311] <= 212;
		weights[312] <= 227;
		weights[313] <= 189;
		weights[314] <= 46;
		weights[315] <= 147;
		weights[316] <= 249;
		weights[317] <= 225;
		weights[318] <= 112;
		weights[319] <= 182;
		weights[320] <= 166;
		weights[321] <= 54;
		weights[322] <= 15;
		weights[323] <= 214;
		weights[324] <= 217;
		weights[325] <= 7;
		weights[326] <= 60;
		weights[327] <= 118;
		weights[328] <= 73;
		weights[329] <= 189;
		weights[330] <= 28;
		weights[331] <= 58;
		weights[332] <= 147;
		weights[333] <= 78;
		weights[334] <= 188;
		weights[335] <= 207;
		weights[336] <= 49;
		weights[337] <= 147;
		weights[338] <= 113;
		weights[339] <= 170;
		weights[340] <= 214;
		weights[341] <= 246;
		weights[342] <= 189;
		weights[343] <= 147;
		weights[344] <= 171;
		weights[345] <= 54;
		weights[346] <= 160;
		weights[347] <= 19;
		weights[348] <= 164;
		weights[349] <= 161;
		weights[350] <= 162;
		weights[351] <= 37;
		weights[352] <= 123;
		weights[353] <= 157;
		weights[354] <= 133;
		weights[355] <= 124;
		weights[356] <= 9;
		weights[357] <= 87;
		weights[358] <= 174;
		weights[359] <= 162;
		weights[360] <= 20;
		weights[361] <= 213;
		weights[362] <= 236;
		weights[363] <= 67;
		weights[364] <= 45;
		weights[365] <= 221;
		weights[366] <= 158;
		weights[367] <= 184;
		weights[368] <= 16;
		weights[369] <= 148;
		weights[370] <= 42;
		weights[371] <= 75;
		weights[372] <= 166;
		weights[373] <= 114;
		weights[374] <= 187;
		weights[375] <= 80;
		weights[376] <= 19;
		weights[377] <= 135;
		weights[378] <= 136;
		weights[379] <= 65;
		weights[380] <= 238;
		weights[381] <= 146;
		weights[382] <= 119;
		weights[383] <= 21;
		weights[384] <= 21;
		weights[385] <= 20;
		weights[386] <= 251;
		weights[387] <= 186;
		weights[388] <= 166;
		weights[389] <= 163;
		weights[390] <= 124;
		weights[391] <= 10;
		weights[392] <= 4;
		weights[393] <= 30;
		weights[394] <= 92;
		weights[395] <= 112;
		weights[396] <= 212;
		weights[397] <= 133;
		weights[398] <= 142;
		weights[399] <= 204;
		weights[400] <= 203;
		weights[401] <= 248;
		weights[402] <= 128;
		weights[403] <= 232;
		weights[404] <= 245;
		weights[405] <= 114;
		weights[406] <= 131;
		weights[407] <= 124;
		weights[408] <= 233;
		weights[409] <= 36;
		weights[410] <= 53;
		weights[411] <= 6;
		weights[412] <= 243;
		weights[413] <= 183;
		weights[414] <= 84;
		weights[415] <= 243;
		weights[416] <= 13;
		weights[417] <= 216;
		weights[418] <= 243;
		weights[419] <= 28;
		weights[420] <= 218;
		weights[421] <= 179;
		weights[422] <= 212;
		weights[423] <= 208;
		weights[424] <= 122;
		weights[425] <= 144;
		weights[426] <= 111;
		weights[427] <= 33;
		weights[428] <= 54;
		weights[429] <= 145;
		weights[430] <= 140;
		weights[431] <= 130;
		weights[432] <= 31;
		weights[433] <= 187;
		weights[434] <= 82;
		weights[435] <= 251;
		weights[436] <= 174;
		weights[437] <= 121;
		weights[438] <= 125;
		weights[439] <= 13;
		weights[440] <= 38;
		weights[441] <= 195;
		weights[442] <= 171;
		weights[443] <= 162;
		weights[444] <= 158;
		weights[445] <= 243;
		weights[446] <= 26;
		weights[447] <= 12;
		weights[448] <= 190;
		weights[449] <= 47;
		weights[450] <= 133;
		weights[451] <= 112;
		weights[452] <= 75;
		weights[453] <= 220;
		weights[454] <= 36;
		weights[455] <= 106;
		weights[456] <= 236;
		weights[457] <= 50;
		weights[458] <= 249;
		weights[459] <= 172;
		weights[460] <= 101;
		weights[461] <= 34;
		weights[462] <= 226;
		weights[463] <= 15;
		weights[464] <= 134;
		weights[465] <= 47;
		weights[466] <= 151;
		weights[467] <= 153;
		weights[468] <= 246;
		weights[469] <= 93;
		weights[470] <= 69;
		weights[471] <= 53;
		weights[472] <= 111;
		weights[473] <= 241;
		weights[474] <= 64;
		weights[475] <= 146;
		weights[476] <= 208;
		weights[477] <= 130;
		weights[478] <= 136;
		weights[479] <= 46;
		weights[480] <= 253;
		weights[481] <= 197;
		weights[482] <= 124;
		weights[483] <= 166;
		weights[484] <= 17;
		weights[485] <= 250;
		weights[486] <= 58;
		weights[487] <= 145;
		weights[488] <= 226;
		weights[489] <= 129;
		weights[490] <= 189;
		weights[491] <= 161;
		weights[492] <= 40;
		weights[493] <= 118;
		weights[494] <= 166;
		weights[495] <= 33;
		weights[496] <= 155;
		weights[497] <= 251;
		weights[498] <= 182;
		weights[499] <= 14;
		weights[500] <= 50;
		weights[501] <= 94;
		weights[502] <= 198;
		weights[503] <= 89;
		weights[504] <= 160;
		weights[505] <= 165;
		weights[506] <= 128;
		weights[507] <= 78;
		weights[508] <= 23;
		weights[509] <= 194;
		weights[510] <= 27;
		weights[511] <= 88;
		weights[512] <= 31;
		weights[513] <= 60;
		weights[514] <= 84;
		weights[515] <= 193;
		weights[516] <= 214;
		weights[517] <= 252;
		weights[518] <= 185;
		weights[519] <= 61;
		weights[520] <= 182;
		weights[521] <= 11;
		weights[522] <= 139;
		weights[523] <= 38;
		weights[524] <= 216;
		weights[525] <= 38;
		weights[526] <= 208;
		weights[527] <= 4;
		weights[528] <= 26;
		weights[529] <= 16;
		weights[530] <= 144;
		weights[531] <= 140;
		weights[532] <= 167;
		weights[533] <= 24;
		weights[534] <= 177;
		weights[535] <= 146;
		weights[536] <= 87;
		weights[537] <= 16;
		weights[538] <= 186;
		weights[539] <= 206;
		weights[540] <= 77;
		weights[541] <= 30;
		weights[542] <= 101;
		weights[543] <= 142;
		weights[544] <= 2;
		weights[545] <= 143;
		weights[546] <= 160;
		weights[547] <= 98;
		weights[548] <= 53;
		weights[549] <= 47;
		weights[550] <= 247;
		weights[551] <= 51;
		weights[552] <= 10;
		weights[553] <= 117;
		weights[554] <= 65;
		weights[555] <= 205;
		weights[556] <= 189;
		weights[557] <= 29;
		weights[558] <= 157;
		weights[559] <= 197;
		weights[560] <= 69;
		weights[561] <= 115;
		weights[562] <= 87;
		weights[563] <= 107;
		weights[564] <= 186;
		weights[565] <= 5;
		weights[566] <= 47;
		weights[567] <= 132;
		weights[568] <= 225;
		weights[569] <= 243;
		weights[570] <= 7;
		weights[571] <= 123;
		weights[572] <= 246;
		weights[573] <= 67;
		weights[574] <= 153;
		weights[575] <= 231;
		weights[576] <= 133;
		weights[577] <= 102;
		weights[578] <= 39;
		weights[579] <= 242;
		weights[580] <= 200;
		weights[581] <= 77;
		weights[582] <= 64;
		weights[583] <= 68;
		weights[584] <= 252;
		weights[585] <= 102;
		weights[586] <= 107;
		weights[587] <= 108;
		weights[588] <= 197;
		weights[589] <= 154;
		weights[590] <= 93;
		weights[591] <= 201;
		weights[592] <= 95;
		weights[593] <= 37;
		weights[594] <= 168;
		weights[595] <= 61;
		weights[596] <= 8;
		weights[597] <= 213;
		weights[598] <= 98;
		weights[599] <= 86;
		weights[600] <= 170;
		weights[601] <= 122;
		weights[602] <= 38;
		weights[603] <= 3;
		weights[604] <= 159;
		weights[605] <= 234;
		weights[606] <= 163;
		weights[607] <= 105;
		weights[608] <= 53;
		weights[609] <= 150;
		weights[610] <= 171;
		weights[611] <= 252;
		weights[612] <= 177;
		weights[613] <= 41;
		weights[614] <= 151;
		weights[615] <= 160;
		weights[616] <= 172;
		weights[617] <= 176;
		weights[618] <= 227;
		weights[619] <= 28;
		weights[620] <= 163;
		weights[621] <= 53;
		weights[622] <= 10;
		weights[623] <= 37;
		weights[624] <= 246;
		weights[625] <= 62;
		weights[626] <= 73;
		weights[627] <= 51;
		weights[628] <= 7;
		weights[629] <= 157;
		weights[630] <= 80;
		weights[631] <= 233;
		weights[632] <= 77;
		weights[633] <= 103;
		weights[634] <= 27;
		weights[635] <= 181;
		weights[636] <= 240;
		weights[637] <= 240;
		weights[638] <= 242;
		weights[639] <= 17;
		weights[640] <= 228;
		weights[641] <= 156;
		weights[642] <= 217;
		weights[643] <= 189;
		weights[644] <= 23;
		weights[645] <= 167;
		weights[646] <= 249;
		weights[647] <= 155;
		weights[648] <= 129;
		weights[649] <= 145;
		weights[650] <= 15;
		weights[651] <= 125;
		weights[652] <= 100;
		weights[653] <= 197;
		weights[654] <= 91;
		weights[655] <= 65;
		weights[656] <= 57;
		weights[657] <= 33;
		weights[658] <= 222;
		weights[659] <= 150;
		weights[660] <= 187;
		weights[661] <= 10;
		weights[662] <= 147;
		weights[663] <= 87;
		weights[664] <= 201;
		weights[665] <= 202;
		weights[666] <= 219;
		weights[667] <= 37;
		weights[668] <= 60;
		weights[669] <= 108;
		weights[670] <= 150;
		weights[671] <= 128;
		weights[672] <= 251;
		weights[673] <= 184;
		weights[674] <= 221;
		weights[675] <= 94;
		weights[676] <= 173;
		weights[677] <= 114;
		weights[678] <= 221;
		weights[679] <= 58;
		weights[680] <= 95;
		weights[681] <= 144;
		weights[682] <= 209;
		weights[683] <= 132;
		weights[684] <= 26;
		weights[685] <= 129;
		weights[686] <= 234;
		weights[687] <= 70;
		weights[688] <= 250;
		weights[689] <= 126;
		weights[690] <= 245;
		weights[691] <= 137;
		weights[692] <= 159;
		weights[693] <= 141;
		weights[694] <= 182;
		weights[695] <= 166;
		weights[696] <= 34;
		weights[697] <= 89;
		weights[698] <= 88;
		weights[699] <= 97;
		weights[700] <= 126;
		weights[701] <= 185;
		weights[702] <= 175;
		weights[703] <= 176;
		weights[704] <= 112;
		weights[705] <= 40;
		weights[706] <= 26;
		weights[707] <= 110;
		weights[708] <= 45;
		weights[709] <= 104;
		weights[710] <= 177;
		weights[711] <= 219;
		weights[712] <= 231;
		weights[713] <= 154;
		weights[714] <= 82;
		weights[715] <= 198;
		weights[716] <= 223;
		weights[717] <= 191;
		weights[718] <= 128;
		weights[719] <= 34;
		weights[720] <= 146;
		weights[721] <= 87;
		weights[722] <= 224;
		weights[723] <= 16;
		weights[724] <= 114;
		weights[725] <= 76;
		weights[726] <= 155;
		weights[727] <= 76;
		weights[728] <= 220;
		weights[729] <= 114;
		weights[730] <= 225;
		weights[731] <= 221;
		weights[732] <= 224;
		weights[733] <= 5;
		weights[734] <= 193;
		weights[735] <= 222;
		weights[736] <= 4;
		weights[737] <= 182;
		weights[738] <= 127;
		weights[739] <= 127;
		weights[740] <= 10;
		weights[741] <= 101;
		weights[742] <= 45;
		weights[743] <= 174;
		weights[744] <= 236;
		weights[745] <= 67;
		weights[746] <= 65;
		weights[747] <= 31;
		weights[748] <= 93;
		weights[749] <= 91;
		weights[750] <= 58;
		weights[751] <= 88;
		weights[752] <= 100;
		weights[753] <= 207;
		weights[754] <= 152;
		weights[755] <= 206;
		weights[756] <= 220;
		weights[757] <= 155;
		weights[758] <= 128;
		weights[759] <= 215;
		weights[760] <= 95;
		weights[761] <= 170;
		weights[762] <= 208;
		weights[763] <= 248;
		weights[764] <= 41;
		weights[765] <= 119;
		weights[766] <= 201;
		weights[767] <= 240;
		weights[768] <= 74;
		weights[769] <= 79;
		weights[770] <= 231;
		weights[771] <= 235;
		weights[772] <= 214;
		weights[773] <= 122;
		weights[774] <= 1;
		weights[775] <= 197;
		weights[776] <= 62;
		weights[777] <= 178;
		weights[778] <= 237;
		weights[779] <= 225;
		weights[780] <= 31;
		weights[781] <= 43;
		weights[782] <= 26;
		weights[783] <= 104;
		weights[784] <= 196;
		weights[785] <= 88;
		weights[786] <= 165;
		weights[787] <= 111;
		weights[788] <= 210;
		weights[789] <= 243;
		weights[790] <= 95;
		weights[791] <= 79;
		weights[792] <= 119;
		weights[793] <= 234;
		weights[794] <= 36;
		weights[795] <= 155;
		weights[796] <= 224;
		weights[797] <= 105;
		weights[798] <= 140;
		weights[799] <= 74;
		weights[800] <= 183;
		weights[801] <= 83;
		weights[802] <= 190;
		weights[803] <= 229;
		weights[804] <= 243;
		weights[805] <= 187;
		weights[806] <= 203;
		weights[807] <= 36;
		weights[808] <= 232;
		weights[809] <= 211;
		weights[810] <= 184;
		weights[811] <= 166;
		weights[812] <= 14;
		weights[813] <= 208;
		weights[814] <= 55;
		weights[815] <= 131;
		weights[816] <= 162;
		weights[817] <= 19;
		weights[818] <= 216;
		weights[819] <= 190;
		weights[820] <= 217;
		weights[821] <= 206;
		weights[822] <= 79;
		weights[823] <= 30;
		weights[824] <= 97;
		weights[825] <= 231;
		weights[826] <= 143;
		weights[827] <= 173;
		weights[828] <= 29;
		weights[829] <= 80;
		weights[830] <= 47;
		weights[831] <= 137;
		weights[832] <= 143;
		weights[833] <= 91;
		weights[834] <= 161;
		weights[835] <= 233;
		weights[836] <= 239;
		weights[837] <= 167;
		weights[838] <= 23;
		weights[839] <= 232;
		weights[840] <= 78;
		weights[841] <= 228;
		weights[842] <= 188;
		weights[843] <= 95;
		weights[844] <= 218;
		weights[845] <= 253;
		weights[846] <= 206;
		weights[847] <= 44;
		weights[848] <= 194;
		weights[849] <= 198;
		weights[850] <= 63;
		weights[851] <= 157;
		weights[852] <= 197;
		weights[853] <= 117;
		weights[854] <= 87;
		weights[855] <= 166;
		weights[856] <= 84;
		weights[857] <= 67;
		weights[858] <= 125;
		weights[859] <= 246;
		weights[860] <= 153;
		weights[861] <= 59;
		weights[862] <= 186;
		weights[863] <= 81;
		weights[864] <= 54;
		weights[865] <= 46;
		weights[866] <= 39;
		weights[867] <= 253;
		weights[868] <= 117;
		weights[869] <= 101;
		weights[870] <= 97;
		weights[871] <= 247;
		weights[872] <= 170;
		weights[873] <= 146;
		weights[874] <= 254;
		weights[875] <= 206;
		weights[876] <= 47;
		weights[877] <= 170;
		weights[878] <= 53;
		weights[879] <= 1;
		weights[880] <= 208;
		weights[881] <= 85;
		weights[882] <= 215;
		weights[883] <= 60;
		weights[884] <= 234;
		weights[885] <= 99;
		weights[886] <= 101;
		weights[887] <= 154;
		weights[888] <= 255;
		weights[889] <= 12;
		weights[890] <= 22;
		weights[891] <= 255;
		weights[892] <= 134;
		weights[893] <= 105;
		weights[894] <= 245;
		weights[895] <= 10;
		weights[896] <= 171;
		weights[897] <= 164;
		weights[898] <= 55;
		weights[899] <= 17;
		weights[900] <= 13;
		weights[901] <= 127;
		weights[902] <= 5;
		weights[903] <= 243;
		weights[904] <= 211;
		weights[905] <= 79;
		weights[906] <= 71;
		weights[907] <= 129;
		weights[908] <= 97;
		weights[909] <= 42;
		weights[910] <= 118;
		weights[911] <= 165;
		weights[912] <= 132;
		weights[913] <= 60;
		weights[914] <= 234;
		weights[915] <= 71;
		weights[916] <= 179;
		weights[917] <= 148;
		weights[918] <= 103;
		weights[919] <= 228;
		weights[920] <= 254;
		weights[921] <= 254;
		weights[922] <= 158;
		weights[923] <= 106;
		weights[924] <= 13;
		weights[925] <= 125;
		weights[926] <= 190;
		weights[927] <= 189;
		weights[928] <= 221;
		weights[929] <= 72;
		weights[930] <= 243;
		weights[931] <= 19;
		weights[932] <= 175;
		weights[933] <= 32;
		weights[934] <= 218;
		weights[935] <= 250;
		weights[936] <= 29;
		weights[937] <= 36;
		weights[938] <= 194;
		weights[939] <= 96;
		weights[940] <= 192;
		weights[941] <= 76;
		weights[942] <= 125;
		weights[943] <= 188;
		weights[944] <= 203;
		weights[945] <= 18;
		weights[946] <= 85;
		weights[947] <= 165;
		weights[948] <= 156;
		weights[949] <= 42;
		weights[950] <= 61;
		weights[951] <= 251;
		weights[952] <= 65;
		weights[953] <= 254;
		weights[954] <= 134;
		weights[955] <= 58;
		weights[956] <= 133;
		weights[957] <= 98;
		weights[958] <= 241;
		weights[959] <= 156;
		weights[960] <= 187;
		weights[961] <= 199;
		weights[962] <= 163;
		weights[963] <= 233;
		weights[964] <= 206;
		weights[965] <= 152;
		weights[966] <= 14;
		weights[967] <= 16;
		weights[968] <= 153;
		weights[969] <= 111;
		weights[970] <= 204;
		weights[971] <= 182;
		weights[972] <= 167;
		weights[973] <= 49;
		weights[974] <= 67;
		weights[975] <= 73;
		weights[976] <= 245;
		weights[977] <= 148;
		weights[978] <= 204;
		weights[979] <= 204;
		weights[980] <= 188;
		weights[981] <= 88;
		weights[982] <= 40;
		weights[983] <= 172;
		weights[984] <= 217;
		weights[985] <= 147;
		weights[986] <= 15;
		weights[987] <= 112;
		weights[988] <= 195;
		weights[989] <= 27;
		weights[990] <= 243;
		weights[991] <= 11;
		weights[992] <= 211;
		weights[993] <= 100;
		weights[994] <= 116;
		weights[995] <= 165;
		weights[996] <= 70;
		weights[997] <= 174;
		weights[998] <= 133;
		weights[999] <= 128;
		weights[1000] <= 85;
		weights[1001] <= 239;
		weights[1002] <= 181;
		weights[1003] <= 90;
		weights[1004] <= 81;
		weights[1005] <= 152;
		weights[1006] <= 11;
		weights[1007] <= 136;
		weights[1008] <= 23;
		weights[1009] <= 94;
		weights[1010] <= 121;
		weights[1011] <= 189;
		weights[1012] <= 166;
		weights[1013] <= 23;
		weights[1014] <= 226;
		weights[1015] <= 203;
		weights[1016] <= 151;
		weights[1017] <= 172;
		weights[1018] <= 244;
		weights[1019] <= 210;
		weights[1020] <= 166;
		weights[1021] <= 157;
		weights[1022] <= 170;
		weights[1023] <= 177;
		weights[1024] <= 218;
		weights[1025] <= 187;
		weights[1026] <= 61;
		weights[1027] <= 112;
		weights[1028] <= 73;
		weights[1029] <= 185;
		weights[1030] <= 11;
		weights[1031] <= 103;
		weights[1032] <= 136;
		weights[1033] <= 3;
		weights[1034] <= 76;
		weights[1035] <= 179;
		weights[1036] <= 183;
		weights[1037] <= 54;
		weights[1038] <= 170;
		weights[1039] <= 134;
		weights[1040] <= 97;
		weights[1041] <= 164;
		weights[1042] <= 14;
		weights[1043] <= 24;
		weights[1044] <= 99;
		weights[1045] <= 113;
		weights[1046] <= 114;
		weights[1047] <= 157;
		weights[1048] <= 162;
		weights[1049] <= 38;
		weights[1050] <= 253;
		weights[1051] <= 179;
		weights[1052] <= 108;
		weights[1053] <= 111;
		weights[1054] <= 160;
		weights[1055] <= 43;
		weights[1056] <= 211;
		weights[1057] <= 19;
		weights[1058] <= 217;
		weights[1059] <= 117;
		weights[1060] <= 37;
		weights[1061] <= 53;
		weights[1062] <= 202;
		weights[1063] <= 11;
		weights[1064] <= 116;
		weights[1065] <= 145;
		weights[1066] <= 209;
		weights[1067] <= 151;
		weights[1068] <= 196;
		weights[1069] <= 64;
		weights[1070] <= 95;
		weights[1071] <= 54;
		weights[1072] <= 124;
		weights[1073] <= 75;
		weights[1074] <= 181;
		weights[1075] <= 100;
		weights[1076] <= 29;
		weights[1077] <= 195;
		weights[1078] <= 55;
		weights[1079] <= 38;
		weights[1080] <= 189;
		weights[1081] <= 17;
		weights[1082] <= 136;
		weights[1083] <= 77;
		weights[1084] <= 90;
		weights[1085] <= 60;
		weights[1086] <= 43;
		weights[1087] <= 81;
		weights[1088] <= 209;
		weights[1089] <= 247;
		weights[1090] <= 225;
		weights[1091] <= 44;
		weights[1092] <= 57;
		weights[1093] <= 86;
		weights[1094] <= 44;
		weights[1095] <= 34;
		weights[1096] <= 193;
		weights[1097] <= 232;
		weights[1098] <= 231;
		weights[1099] <= 122;
		weights[1100] <= 236;
		weights[1101] <= 179;
		weights[1102] <= 166;
		weights[1103] <= 214;
		weights[1104] <= 223;
		weights[1105] <= 65;
		weights[1106] <= 64;
		weights[1107] <= 192;
		weights[1108] <= 30;
		weights[1109] <= 160;
		weights[1110] <= 44;
		weights[1111] <= 215;
		weights[1112] <= 99;
		weights[1113] <= 52;
		weights[1114] <= 148;
		weights[1115] <= 234;
		weights[1116] <= 44;
		weights[1117] <= 234;
		weights[1118] <= 105;
		weights[1119] <= 229;
		weights[1120] <= 248;
		weights[1121] <= 152;
		weights[1122] <= 42;
		weights[1123] <= 209;
		weights[1124] <= 241;
		weights[1125] <= 212;
		weights[1126] <= 246;
		weights[1127] <= 22;
		weights[1128] <= 32;
		weights[1129] <= 98;
		weights[1130] <= 26;
		weights[1131] <= 140;
		weights[1132] <= 22;
		weights[1133] <= 248;
		weights[1134] <= 171;
		weights[1135] <= 88;
		weights[1136] <= 62;
		weights[1137] <= 251;
		weights[1138] <= 210;
		weights[1139] <= 22;
		weights[1140] <= 72;
		weights[1141] <= 102;
		weights[1142] <= 60;
		weights[1143] <= 34;
		weights[1144] <= 10;
		weights[1145] <= 132;
		weights[1146] <= 113;
		weights[1147] <= 165;
		weights[1148] <= 150;
		weights[1149] <= 247;
		weights[1150] <= 224;
		weights[1151] <= 93;
		weights[1152] <= 241;
		weights[1153] <= 48;
		weights[1154] <= 70;
		weights[1155] <= 97;
		weights[1156] <= 80;
		weights[1157] <= 194;
		weights[1158] <= 174;
		weights[1159] <= 64;
		weights[1160] <= 245;
		weights[1161] <= 244;
		weights[1162] <= 228;
		weights[1163] <= 61;
		weights[1164] <= 33;
		weights[1165] <= 112;
		weights[1166] <= 24;
		weights[1167] <= 221;
		weights[1168] <= 167;
		weights[1169] <= 59;
		weights[1170] <= 126;
		weights[1171] <= 196;
		weights[1172] <= 61;
		weights[1173] <= 137;
		weights[1174] <= 136;
		weights[1175] <= 213;
		weights[1176] <= 25;
		weights[1177] <= 19;
		weights[1178] <= 23;
		weights[1179] <= 58;
		weights[1180] <= 249;
		weights[1181] <= 100;
		weights[1182] <= 173;
		weights[1183] <= 134;
		weights[1184] <= 161;
		weights[1185] <= 153;
		weights[1186] <= 233;
		weights[1187] <= 42;
		weights[1188] <= 97;
		weights[1189] <= 197;
		weights[1190] <= 134;
		weights[1191] <= 138;
		weights[1192] <= 216;
		weights[1193] <= 199;
		weights[1194] <= 26;
		weights[1195] <= 90;
		weights[1196] <= 78;
		weights[1197] <= 177;
		weights[1198] <= 128;
		weights[1199] <= 74;
		weights[1200] <= 24;
		weights[1201] <= 10;
		weights[1202] <= 180;
		weights[1203] <= 31;
		weights[1204] <= 30;
		weights[1205] <= 173;
		weights[1206] <= 188;
		weights[1207] <= 184;
		weights[1208] <= 166;
		weights[1209] <= 56;
		weights[1210] <= 35;
		weights[1211] <= 145;
		weights[1212] <= 20;
		weights[1213] <= 14;
		weights[1214] <= 218;
		weights[1215] <= 240;
		weights[1216] <= 157;
		weights[1217] <= 102;
		weights[1218] <= 19;
		weights[1219] <= 34;
		weights[1220] <= 160;
		weights[1221] <= 53;
		weights[1222] <= 161;
		weights[1223] <= 23;
		weights[1224] <= 155;
		weights[1225] <= 218;
		weights[1226] <= 230;
		weights[1227] <= 240;
		weights[1228] <= 241;
		weights[1229] <= 62;
		weights[1230] <= 242;
		weights[1231] <= 223;
		weights[1232] <= 154;
		weights[1233] <= 96;
		weights[1234] <= 224;
		weights[1235] <= 187;
		weights[1236] <= 91;
		weights[1237] <= 246;
		weights[1238] <= 70;
		weights[1239] <= 159;
		weights[1240] <= 147;
		weights[1241] <= 128;
		weights[1242] <= 155;
		weights[1243] <= 53;
		weights[1244] <= 106;
		weights[1245] <= 24;
		weights[1246] <= 198;
		weights[1247] <= 109;
		weights[1248] <= 130;
		weights[1249] <= 101;
		weights[1250] <= 119;
		weights[1251] <= 148;
		weights[1252] <= 219;
		weights[1253] <= 218;
		weights[1254] <= 101;
		weights[1255] <= 72;
		weights[1256] <= 180;
		weights[1257] <= 141;
		weights[1258] <= 207;
		weights[1259] <= 84;
		weights[1260] <= 61;
		weights[1261] <= 239;
		weights[1262] <= 159;
		weights[1263] <= 143;
		weights[1264] <= 162;
		weights[1265] <= 80;
		weights[1266] <= 192;
		weights[1267] <= 203;
		weights[1268] <= 105;
		weights[1269] <= 225;
		weights[1270] <= 76;
		weights[1271] <= 7;
		weights[1272] <= 254;
		weights[1273] <= 243;
		weights[1274] <= 28;
		weights[1275] <= 138;
		weights[1276] <= 167;
		weights[1277] <= 187;
		weights[1278] <= 8;
		weights[1279] <= 27;
		weights[1280] <= 30;
		weights[1281] <= 249;
		weights[1282] <= 83;
		weights[1283] <= 34;
		weights[1284] <= 24;
		weights[1285] <= 107;
		weights[1286] <= 168;
		weights[1287] <= 121;
		weights[1288] <= 48;
		weights[1289] <= 144;
		weights[1290] <= 145;
		weights[1291] <= 13;
		weights[1292] <= 121;
		weights[1293] <= 3;
		weights[1294] <= 248;
		weights[1295] <= 134;
		weights[1296] <= 118;
		weights[1297] <= 179;
		weights[1298] <= 25;
		weights[1299] <= 88;
		weights[1300] <= 176;
		weights[1301] <= 242;
		weights[1302] <= 177;
		weights[1303] <= 229;
		weights[1304] <= 243;
		weights[1305] <= 199;
		weights[1306] <= 58;
		weights[1307] <= 44;
		weights[1308] <= 63;
		weights[1309] <= 12;
		weights[1310] <= 137;
		weights[1311] <= 203;
		weights[1312] <= 143;
		weights[1313] <= 89;
		weights[1314] <= 137;
		weights[1315] <= 250;
		weights[1316] <= 215;
		weights[1317] <= 197;
		weights[1318] <= 232;
		weights[1319] <= 24;
		weights[1320] <= 88;
		weights[1321] <= 244;
		weights[1322] <= 49;
		weights[1323] <= 117;
		weights[1324] <= 136;
		weights[1325] <= 147;
		weights[1326] <= 153;
		weights[1327] <= 161;
		weights[1328] <= 75;
		weights[1329] <= 173;
		weights[1330] <= 255;
		weights[1331] <= 20;
		weights[1332] <= 94;
		weights[1333] <= 111;
		weights[1334] <= 74;
		weights[1335] <= 97;
		weights[1336] <= 201;
		weights[1337] <= 53;
		weights[1338] <= 111;
		weights[1339] <= 171;
		weights[1340] <= 12;
		weights[1341] <= 20;
		weights[1342] <= 238;
		weights[1343] <= 27;
		weights[1344] <= 12;
		weights[1345] <= 168;
		weights[1346] <= 3;
		weights[1347] <= 182;
		weights[1348] <= 62;
		weights[1349] <= 241;
		weights[1350] <= 103;
		weights[1351] <= 52;
		weights[1352] <= 161;
		weights[1353] <= 190;
		weights[1354] <= 98;
		weights[1355] <= 46;
		weights[1356] <= 149;
		weights[1357] <= 87;
		weights[1358] <= 42;
		weights[1359] <= 96;
		weights[1360] <= 104;
		weights[1361] <= 212;
		weights[1362] <= 233;
		weights[1363] <= 31;
		weights[1364] <= 27;
		weights[1365] <= 171;
		weights[1366] <= 43;
		weights[1367] <= 87;
		weights[1368] <= 79;
		weights[1369] <= 163;
		weights[1370] <= 114;
		weights[1371] <= 146;
		weights[1372] <= 91;
		weights[1373] <= 190;
		weights[1374] <= 102;
		weights[1375] <= 165;
		weights[1376] <= 106;
		weights[1377] <= 234;
		weights[1378] <= 116;
		weights[1379] <= 20;
		weights[1380] <= 218;
		weights[1381] <= 240;
		weights[1382] <= 48;
		weights[1383] <= 237;
		weights[1384] <= 117;
		weights[1385] <= 59;
		weights[1386] <= 215;
		weights[1387] <= 203;
		weights[1388] <= 32;
		weights[1389] <= 220;
		weights[1390] <= 171;
		weights[1391] <= 218;
		weights[1392] <= 239;
		weights[1393] <= 195;
		weights[1394] <= 195;
		weights[1395] <= 193;
		weights[1396] <= 133;
		weights[1397] <= 216;
		weights[1398] <= 2;
		weights[1399] <= 204;
		weights[1400] <= 87;
		weights[1401] <= 143;
		weights[1402] <= 168;
		weights[1403] <= 23;
		weights[1404] <= 137;
		weights[1405] <= 215;
		weights[1406] <= 142;
		weights[1407] <= 109;
		weights[1408] <= 184;
		weights[1409] <= 99;
		weights[1410] <= 170;
		weights[1411] <= 124;
		weights[1412] <= 143;
		weights[1413] <= 174;
		weights[1414] <= 192;
		weights[1415] <= 14;
		weights[1416] <= 52;
		weights[1417] <= 15;
		weights[1418] <= 123;
		weights[1419] <= 47;
		weights[1420] <= 19;
		weights[1421] <= 225;
		weights[1422] <= 179;
		weights[1423] <= 137;
		weights[1424] <= 143;
		weights[1425] <= 238;
		weights[1426] <= 163;
		weights[1427] <= 104;
		weights[1428] <= 8;
		weights[1429] <= 226;
		weights[1430] <= 167;
		weights[1431] <= 17;
		weights[1432] <= 125;
		weights[1433] <= 175;
		weights[1434] <= 239;
		weights[1435] <= 160;
		weights[1436] <= 45;
		weights[1437] <= 114;
		weights[1438] <= 24;
		weights[1439] <= 159;
		weights[1440] <= 254;
		weights[1441] <= 89;
		weights[1442] <= 131;
		weights[1443] <= 179;
		weights[1444] <= 95;
		weights[1445] <= 234;
		weights[1446] <= 103;
		weights[1447] <= 253;
		weights[1448] <= 195;
		weights[1449] <= 130;
		weights[1450] <= 178;
		weights[1451] <= 204;
		weights[1452] <= 244;
		weights[1453] <= 194;
		weights[1454] <= 26;
		weights[1455] <= 153;
		weights[1456] <= 138;
		weights[1457] <= 163;
		weights[1458] <= 33;
		weights[1459] <= 216;
		weights[1460] <= 98;
		weights[1461] <= 123;
		weights[1462] <= 249;
		weights[1463] <= 94;
		weights[1464] <= 208;
		weights[1465] <= 105;
		weights[1466] <= 249;
		weights[1467] <= 40;
		weights[1468] <= 94;
		weights[1469] <= 188;
		weights[1470] <= 239;
		weights[1471] <= 93;
		weights[1472] <= 169;
		weights[1473] <= 27;
		weights[1474] <= 179;
		weights[1475] <= 204;
		weights[1476] <= 90;
		weights[1477] <= 208;
		weights[1478] <= 181;
		weights[1479] <= 40;
		weights[1480] <= 45;
		weights[1481] <= 208;
		weights[1482] <= 211;
		weights[1483] <= 211;
		weights[1484] <= 161;
		weights[1485] <= 255;
		weights[1486] <= 9;
		weights[1487] <= 22;
		weights[1488] <= 164;
		weights[1489] <= 55;
		weights[1490] <= 60;
		weights[1491] <= 38;
		weights[1492] <= 191;
		weights[1493] <= 242;
		weights[1494] <= 121;
		weights[1495] <= 243;
		weights[1496] <= 248;
		weights[1497] <= 137;
		weights[1498] <= 28;
		weights[1499] <= 251;
		weights[1500] <= 238;
		weights[1501] <= 77;
		weights[1502] <= 234;
		weights[1503] <= 94;
		weights[1504] <= 178;
		weights[1505] <= 219;
		weights[1506] <= 99;
		weights[1507] <= 53;
		weights[1508] <= 126;
		weights[1509] <= 110;
		weights[1510] <= 20;
		weights[1511] <= 139;
		weights[1512] <= 62;
		weights[1513] <= 253;
		weights[1514] <= 227;
		weights[1515] <= 195;
		weights[1516] <= 20;
		weights[1517] <= 233;
		weights[1518] <= 97;
		weights[1519] <= 196;
		weights[1520] <= 82;
		weights[1521] <= 22;
		weights[1522] <= 244;
		weights[1523] <= 124;
		weights[1524] <= 34;
		weights[1525] <= 182;
		weights[1526] <= 246;
		weights[1527] <= 140;
		weights[1528] <= 251;
		weights[1529] <= 11;
		weights[1530] <= 109;
		weights[1531] <= 143;
		weights[1532] <= 86;
		weights[1533] <= 105;
		weights[1534] <= 90;
		weights[1535] <= 103;
		weights[1536] <= 6;
		weights[1537] <= 222;
		weights[1538] <= 146;
		weights[1539] <= 120;
		weights[1540] <= 88;
		weights[1541] <= 60;
		weights[1542] <= 117;
		weights[1543] <= 210;
		weights[1544] <= 5;
		weights[1545] <= 245;
		weights[1546] <= 51;
		weights[1547] <= 178;
		weights[1548] <= 30;
		weights[1549] <= 185;
		weights[1550] <= 197;
		weights[1551] <= 14;
		weights[1552] <= 81;
		weights[1553] <= 26;
		weights[1554] <= 70;
		weights[1555] <= 211;
		weights[1556] <= 227;
		weights[1557] <= 122;
		weights[1558] <= 205;
		weights[1559] <= 186;
		weights[1560] <= 107;
		weights[1561] <= 168;
		weights[1562] <= 237;
		weights[1563] <= 64;
		weights[1564] <= 38;
		weights[1565] <= 142;
		weights[1566] <= 101;
		weights[1567] <= 204;
		weights[1568] <= 6;
		weights[1569] <= 227;
		weights[1570] <= 45;
		weights[1571] <= 17;
		weights[1572] <= 50;
		weights[1573] <= 171;
		weights[1574] <= 243;
		weights[1575] <= 66;
		weights[1576] <= 198;
		weights[1577] <= 145;
		weights[1578] <= 68;
		weights[1579] <= 153;
		weights[1580] <= 186;
		weights[1581] <= 19;
		weights[1582] <= 210;
		weights[1583] <= 231;
		weights[1584] <= 229;
		weights[1585] <= 123;
		weights[1586] <= 97;
		weights[1587] <= 237;
		weights[1588] <= 115;
		weights[1589] <= 178;
		weights[1590] <= 33;
		weights[1591] <= 91;
		weights[1592] <= 167;
		weights[1593] <= 52;
		weights[1594] <= 62;
		weights[1595] <= 110;
		weights[1596] <= 81;
		weights[1597] <= 188;
		weights[1598] <= 229;
		weights[1599] <= 127;
		weights[1600] <= 219;
		weights[1601] <= 176;
		weights[1602] <= 90;
		weights[1603] <= 255;
		weights[1604] <= 37;
		weights[1605] <= 237;
		weights[1606] <= 29;
		weights[1607] <= 42;
		weights[1608] <= 92;
		weights[1609] <= 170;
		weights[1610] <= 192;
		weights[1611] <= 75;
		weights[1612] <= 108;
		weights[1613] <= 223;
		weights[1614] <= 113;
		weights[1615] <= 95;
		weights[1616] <= 77;
		weights[1617] <= 146;
		weights[1618] <= 80;
		weights[1619] <= 138;
		weights[1620] <= 194;
		weights[1621] <= 103;
		weights[1622] <= 201;
		weights[1623] <= 237;
		weights[1624] <= 179;
		weights[1625] <= 19;
		weights[1626] <= 101;
		weights[1627] <= 75;
		weights[1628] <= 114;
		weights[1629] <= 6;
		weights[1630] <= 227;
		weights[1631] <= 134;
		weights[1632] <= 226;
		weights[1633] <= 252;
		weights[1634] <= 188;
		weights[1635] <= 135;
		weights[1636] <= 48;
		weights[1637] <= 202;
		weights[1638] <= 82;
		weights[1639] <= 228;
		weights[1640] <= 11;
		weights[1641] <= 246;
		weights[1642] <= 247;
		weights[1643] <= 123;
		weights[1644] <= 208;
		weights[1645] <= 240;
		weights[1646] <= 37;
		weights[1647] <= 154;
		weights[1648] <= 66;
		weights[1649] <= 12;
		weights[1650] <= 25;
		weights[1651] <= 216;
		weights[1652] <= 82;
		weights[1653] <= 60;
		weights[1654] <= 131;
		weights[1655] <= 47;
		weights[1656] <= 109;
		weights[1657] <= 32;
		weights[1658] <= 34;
		weights[1659] <= 65;
		weights[1660] <= 117;
		weights[1661] <= 214;
		weights[1662] <= 196;
		weights[1663] <= 33;
		weights[1664] <= 57;
		weights[1665] <= 8;
		weights[1666] <= 172;
		weights[1667] <= 148;
		weights[1668] <= 190;
		weights[1669] <= 121;
		weights[1670] <= 118;
		weights[1671] <= 242;
		weights[1672] <= 167;
		weights[1673] <= 116;
		weights[1674] <= 227;
		weights[1675] <= 111;
		weights[1676] <= 163;
		weights[1677] <= 18;
		weights[1678] <= 241;
		weights[1679] <= 164;
		weights[1680] <= 175;
		weights[1681] <= 42;
		weights[1682] <= 62;
		weights[1683] <= 8;
		weights[1684] <= 136;
		weights[1685] <= 138;
		weights[1686] <= 7;
		weights[1687] <= 93;
		weights[1688] <= 228;
		weights[1689] <= 184;
		weights[1690] <= 27;
		weights[1691] <= 37;
		weights[1692] <= 179;
		weights[1693] <= 91;
		weights[1694] <= 175;
		weights[1695] <= 25;
		weights[1696] <= 119;
		weights[1697] <= 164;
		weights[1698] <= 217;
		weights[1699] <= 236;
		weights[1700] <= 55;
		weights[1701] <= 208;
		weights[1702] <= 198;
		weights[1703] <= 185;
		weights[1704] <= 233;
		weights[1705] <= 205;
		weights[1706] <= 247;
		weights[1707] <= 134;
		weights[1708] <= 213;
		weights[1709] <= 108;
		weights[1710] <= 74;
		weights[1711] <= 206;
		weights[1712] <= 137;
		weights[1713] <= 215;
		weights[1714] <= 110;
		weights[1715] <= 170;
		weights[1716] <= 178;
		weights[1717] <= 191;
		weights[1718] <= 136;
		weights[1719] <= 134;
		weights[1720] <= 224;
		weights[1721] <= 21;
		weights[1722] <= 113;
		weights[1723] <= 112;
		weights[1724] <= 35;
		weights[1725] <= 69;
		weights[1726] <= 40;
		weights[1727] <= 223;
		weights[1728] <= 31;
		weights[1729] <= 221;
		weights[1730] <= 141;
		weights[1731] <= 219;
		weights[1732] <= 138;
		weights[1733] <= 20;
		weights[1734] <= 61;
		weights[1735] <= 50;
		weights[1736] <= 220;
		weights[1737] <= 82;
		weights[1738] <= 76;
		weights[1739] <= 255;
		weights[1740] <= 122;
		weights[1741] <= 115;
		weights[1742] <= 162;
		weights[1743] <= 255;
		weights[1744] <= 59;
		weights[1745] <= 93;
		weights[1746] <= 88;
		weights[1747] <= 40;
		weights[1748] <= 112;
		weights[1749] <= 140;
		weights[1750] <= 184;
		weights[1751] <= 82;
		weights[1752] <= 68;
		weights[1753] <= 180;
		weights[1754] <= 38;
		weights[1755] <= 118;
		weights[1756] <= 196;
		weights[1757] <= 183;
		weights[1758] <= 45;
		weights[1759] <= 97;
		weights[1760] <= 147;
		weights[1761] <= 213;
		weights[1762] <= 224;
		weights[1763] <= 78;
		weights[1764] <= 44;
		weights[1765] <= 84;
		weights[1766] <= 92;
		weights[1767] <= 221;
		weights[1768] <= 119;
		weights[1769] <= 155;
		weights[1770] <= 57;
		weights[1771] <= 115;
		weights[1772] <= 99;
		weights[1773] <= 138;
		weights[1774] <= 186;
		weights[1775] <= 78;
		weights[1776] <= 188;
		weights[1777] <= 77;
		weights[1778] <= 123;
		weights[1779] <= 93;
		weights[1780] <= 206;
		weights[1781] <= 58;
		weights[1782] <= 17;
		weights[1783] <= 94;
		weights[1784] <= 174;
		weights[1785] <= 228;
		weights[1786] <= 17;
		weights[1787] <= 9;
		weights[1788] <= 182;
		weights[1789] <= 54;
		weights[1790] <= 189;
		weights[1791] <= 61;
		weights[1792] <= 166;
		weights[1793] <= 53;
		weights[1794] <= 169;
		weights[1795] <= 73;
		weights[1796] <= 209;
		weights[1797] <= 95;
		weights[1798] <= 95;
		weights[1799] <= 252;
		weights[1800] <= 251;
		weights[1801] <= 62;
		weights[1802] <= 233;
		weights[1803] <= 32;
		weights[1804] <= 219;
		weights[1805] <= 157;
		weights[1806] <= 203;
		weights[1807] <= 28;
		weights[1808] <= 79;
		weights[1809] <= 240;
		weights[1810] <= 255;
		weights[1811] <= 103;
		weights[1812] <= 27;
		weights[1813] <= 117;
		weights[1814] <= 83;
		weights[1815] <= 88;
		weights[1816] <= 174;
		weights[1817] <= 255;
		weights[1818] <= 96;
		weights[1819] <= 222;
		weights[1820] <= 67;
		weights[1821] <= 165;
		weights[1822] <= 222;
		weights[1823] <= 182;
		weights[1824] <= 27;
		weights[1825] <= 191;
		weights[1826] <= 82;
		weights[1827] <= 91;
		weights[1828] <= 157;
		weights[1829] <= 156;
		weights[1830] <= 249;
		weights[1831] <= 128;
		weights[1832] <= 71;
		weights[1833] <= 25;
		weights[1834] <= 209;
		weights[1835] <= 78;
		weights[1836] <= 8;
		weights[1837] <= 104;
		weights[1838] <= 3;
		weights[1839] <= 252;
		weights[1840] <= 205;
		weights[1841] <= 44;
		weights[1842] <= 109;
		weights[1843] <= 161;
		weights[1844] <= 143;
		weights[1845] <= 29;
		weights[1846] <= 180;
		weights[1847] <= 28;
		weights[1848] <= 63;
		weights[1849] <= 148;
		weights[1850] <= 186;
		weights[1851] <= 217;
		weights[1852] <= 246;
		weights[1853] <= 243;
		weights[1854] <= 77;
		weights[1855] <= 97;
		weights[1856] <= 246;
		weights[1857] <= 194;
		weights[1858] <= 111;
		weights[1859] <= 162;
		weights[1860] <= 10;
		weights[1861] <= 159;
		weights[1862] <= 129;
		weights[1863] <= 144;
		weights[1864] <= 75;
		weights[1865] <= 224;
		weights[1866] <= 247;
		weights[1867] <= 88;
		weights[1868] <= 64;
		weights[1869] <= 24;
		weights[1870] <= 189;
		weights[1871] <= 78;
		weights[1872] <= 72;
		weights[1873] <= 212;
		weights[1874] <= 196;
		weights[1875] <= 72;
		weights[1876] <= 171;
		weights[1877] <= 234;
		weights[1878] <= 72;
		weights[1879] <= 58;
		weights[1880] <= 185;
		weights[1881] <= 159;
		weights[1882] <= 26;
		weights[1883] <= 32;
		weights[1884] <= 35;
		weights[1885] <= 45;
		weights[1886] <= 89;
		weights[1887] <= 122;
		weights[1888] <= 116;
		weights[1889] <= 165;
		weights[1890] <= 147;
		weights[1891] <= 195;
		weights[1892] <= 36;
		weights[1893] <= 120;
		weights[1894] <= 208;
		weights[1895] <= 40;
		weights[1896] <= 75;
		weights[1897] <= 14;
		weights[1898] <= 150;
		weights[1899] <= 198;
		weights[1900] <= 29;
		weights[1901] <= 188;
		weights[1902] <= 218;
		weights[1903] <= 136;
		weights[1904] <= 148;
		weights[1905] <= 3;
		weights[1906] <= 69;
		weights[1907] <= 191;
		weights[1908] <= 145;
		weights[1909] <= 234;
		weights[1910] <= 71;
		weights[1911] <= 3;
		weights[1912] <= 49;
		weights[1913] <= 54;
		weights[1914] <= 193;
		weights[1915] <= 20;
		weights[1916] <= 93;
		weights[1917] <= 15;
		weights[1918] <= 228;
		weights[1919] <= 23;
		weights[1920] <= 22;
		weights[1921] <= 195;
		weights[1922] <= 133;
		weights[1923] <= 87;
		weights[1924] <= 236;
		weights[1925] <= 94;
		weights[1926] <= 196;
		weights[1927] <= 149;
		weights[1928] <= 191;
		weights[1929] <= 241;
		weights[1930] <= 54;
		weights[1931] <= 28;
		weights[1932] <= 132;
		weights[1933] <= 74;
		weights[1934] <= 91;
		weights[1935] <= 11;
		weights[1936] <= 239;
		weights[1937] <= 68;
		weights[1938] <= 92;
		weights[1939] <= 214;
		weights[1940] <= 2;
		weights[1941] <= 221;
		weights[1942] <= 95;
		weights[1943] <= 80;
		weights[1944] <= 48;
		weights[1945] <= 120;
		weights[1946] <= 207;
		weights[1947] <= 64;
		weights[1948] <= 193;
		weights[1949] <= 130;
		weights[1950] <= 234;
		weights[1951] <= 27;
		weights[1952] <= 211;
		weights[1953] <= 7;
		weights[1954] <= 48;
		weights[1955] <= 136;
		weights[1956] <= 78;
		weights[1957] <= 96;
		weights[1958] <= 104;
		weights[1959] <= 7;
		weights[1960] <= 151;
		weights[1961] <= 95;
		weights[1962] <= 153;
		weights[1963] <= 175;
		weights[1964] <= 14;
		weights[1965] <= 255;
		weights[1966] <= 41;
		weights[1967] <= 77;
		weights[1968] <= 160;
		weights[1969] <= 9;
		weights[1970] <= 193;
		weights[1971] <= 170;
		weights[1972] <= 89;
		weights[1973] <= 39;
		weights[1974] <= 146;
		weights[1975] <= 236;
		weights[1976] <= 102;
		weights[1977] <= 217;
		weights[1978] <= 130;
		weights[1979] <= 98;
		weights[1980] <= 171;
		weights[1981] <= 161;
		weights[1982] <= 29;
		weights[1983] <= 116;
		weights[1984] <= 127;
		weights[1985] <= 63;
		weights[1986] <= 21;
		weights[1987] <= 186;
		weights[1988] <= 217;
		weights[1989] <= 16;
		weights[1990] <= 191;
		weights[1991] <= 15;
		weights[1992] <= 74;
		weights[1993] <= 166;
		weights[1994] <= 124;
		weights[1995] <= 162;
		weights[1996] <= 7;
		weights[1997] <= 188;
		weights[1998] <= 224;
		weights[1999] <= 158;
		weights[2000] <= 152;
		weights[2001] <= 66;
		weights[2002] <= 160;
		weights[2003] <= 243;
		weights[2004] <= 217;
		weights[2005] <= 196;
		weights[2006] <= 139;
		weights[2007] <= 245;
		weights[2008] <= 147;
		weights[2009] <= 215;
		weights[2010] <= 218;
		weights[2011] <= 126;
		weights[2012] <= 176;
		weights[2013] <= 13;
		weights[2014] <= 244;
		weights[2015] <= 218;
		weights[2016] <= 201;
		weights[2017] <= 185;
		weights[2018] <= 215;
		weights[2019] <= 100;
		weights[2020] <= 57;
		weights[2021] <= 233;
		weights[2022] <= 197;
		weights[2023] <= 89;
		weights[2024] <= 189;
		weights[2025] <= 65;
		weights[2026] <= 28;
		weights[2027] <= 222;
		weights[2028] <= 145;
		weights[2029] <= 172;
		weights[2030] <= 105;
		weights[2031] <= 191;
		weights[2032] <= 232;
		weights[2033] <= 88;
		weights[2034] <= 219;
		weights[2035] <= 26;
		weights[2036] <= 152;
		weights[2037] <= 145;
		weights[2038] <= 5;
		weights[2039] <= 62;
		weights[2040] <= 154;
		weights[2041] <= 96;
		weights[2042] <= 206;
		weights[2043] <= 145;
		weights[2044] <= 243;
		weights[2045] <= 9;
		weights[2046] <= 197;
		weights[2047] <= 187;
		weights[2048] <= 111;
		weights[2049] <= 230;
		weights[2050] <= 213;
		weights[2051] <= 154;
		weights[2052] <= 46;
		weights[2053] <= 143;
		weights[2054] <= 121;
		weights[2055] <= 224;
		weights[2056] <= 79;
		weights[2057] <= 219;
		weights[2058] <= 228;
		weights[2059] <= 128;
		weights[2060] <= 142;
		weights[2061] <= 38;
		weights[2062] <= 186;
		weights[2063] <= 232;
		weights[2064] <= 246;
		weights[2065] <= 7;
		weights[2066] <= 50;
		weights[2067] <= 17;
		weights[2068] <= 22;
		weights[2069] <= 27;
		weights[2070] <= 97;
		weights[2071] <= 19;
		weights[2072] <= 167;
		weights[2073] <= 85;
		weights[2074] <= 238;
		weights[2075] <= 191;
		weights[2076] <= 149;
		weights[2077] <= 58;
		weights[2078] <= 107;
		weights[2079] <= 2;
		weights[2080] <= 187;
		weights[2081] <= 19;
		weights[2082] <= 15;
		weights[2083] <= 31;
		weights[2084] <= 225;
		weights[2085] <= 58;
		weights[2086] <= 49;
		weights[2087] <= 187;
		weights[2088] <= 198;
		weights[2089] <= 84;
		weights[2090] <= 213;
		weights[2091] <= 140;
		weights[2092] <= 180;
		weights[2093] <= 108;
		weights[2094] <= 116;
		weights[2095] <= 114;
		weights[2096] <= 223;
		weights[2097] <= 119;
		weights[2098] <= 138;
		weights[2099] <= 55;
		weights[2100] <= 196;
		weights[2101] <= 193;
		weights[2102] <= 194;
		weights[2103] <= 106;
		weights[2104] <= 38;
		weights[2105] <= 239;
		weights[2106] <= 246;
		weights[2107] <= 91;
		weights[2108] <= 37;
		weights[2109] <= 2;
		weights[2110] <= 28;
		weights[2111] <= 12;
		weights[2112] <= 42;
		weights[2113] <= 102;
		weights[2114] <= 155;
		weights[2115] <= 36;
		weights[2116] <= 216;
		weights[2117] <= 3;
		weights[2118] <= 67;
		weights[2119] <= 33;
		weights[2120] <= 134;
		weights[2121] <= 26;
		weights[2122] <= 192;
		weights[2123] <= 161;
		weights[2124] <= 66;
		weights[2125] <= 138;
		weights[2126] <= 140;
		weights[2127] <= 194;
		weights[2128] <= 136;
		weights[2129] <= 2;
		weights[2130] <= 17;
		weights[2131] <= 24;
		weights[2132] <= 111;
		weights[2133] <= 39;
		weights[2134] <= 124;
		weights[2135] <= 240;
		weights[2136] <= 164;
		weights[2137] <= 238;
		weights[2138] <= 198;
		weights[2139] <= 131;
		weights[2140] <= 17;
		weights[2141] <= 76;
		weights[2142] <= 17;
		weights[2143] <= 79;
		weights[2144] <= 211;
		weights[2145] <= 35;
		weights[2146] <= 135;
		weights[2147] <= 180;
		weights[2148] <= 253;
		weights[2149] <= 142;
		weights[2150] <= 33;
		weights[2151] <= 149;
		weights[2152] <= 159;
		weights[2153] <= 162;
		weights[2154] <= 168;
		weights[2155] <= 81;
		weights[2156] <= 244;
		weights[2157] <= 243;
		weights[2158] <= 43;
		weights[2159] <= 7;
		weights[2160] <= 21;
		weights[2161] <= 209;
		weights[2162] <= 93;
		weights[2163] <= 220;
		weights[2164] <= 16;
		weights[2165] <= 81;
		weights[2166] <= 25;
		weights[2167] <= 160;
		weights[2168] <= 34;
		weights[2169] <= 31;
		weights[2170] <= 61;
		weights[2171] <= 243;
		weights[2172] <= 172;
		weights[2173] <= 179;
		weights[2174] <= 88;
		weights[2175] <= 251;
		weights[2176] <= 22;
		weights[2177] <= 255;
		weights[2178] <= 141;
		weights[2179] <= 188;
		weights[2180] <= 23;
		weights[2181] <= 116;
		weights[2182] <= 252;
		weights[2183] <= 216;
		weights[2184] <= 231;
		weights[2185] <= 51;
		weights[2186] <= 67;
		weights[2187] <= 69;
		weights[2188] <= 249;
		weights[2189] <= 58;
		weights[2190] <= 25;
		weights[2191] <= 179;
		weights[2192] <= 169;
		weights[2193] <= 178;
		weights[2194] <= 201;
		weights[2195] <= 107;
		weights[2196] <= 133;
		weights[2197] <= 167;
		weights[2198] <= 197;
		weights[2199] <= 101;
		weights[2200] <= 31;
		weights[2201] <= 179;
		weights[2202] <= 38;
		weights[2203] <= 160;
		weights[2204] <= 23;
		weights[2205] <= 35;
		weights[2206] <= 181;
		weights[2207] <= 190;
		weights[2208] <= 72;
		weights[2209] <= 5;
		weights[2210] <= 121;
		weights[2211] <= 131;
		weights[2212] <= 40;
		weights[2213] <= 71;
		weights[2214] <= 211;
		weights[2215] <= 173;
		weights[2216] <= 100;
		weights[2217] <= 70;
		weights[2218] <= 240;
		weights[2219] <= 74;
		weights[2220] <= 141;
		weights[2221] <= 119;
		weights[2222] <= 106;
		weights[2223] <= 65;
		weights[2224] <= 236;
		weights[2225] <= 206;
		weights[2226] <= 47;
		weights[2227] <= 159;
		weights[2228] <= 70;
		weights[2229] <= 56;
		weights[2230] <= 231;
		weights[2231] <= 250;
		weights[2232] <= 116;
		weights[2233] <= 98;
		weights[2234] <= 44;
		weights[2235] <= 226;
		weights[2236] <= 73;
		weights[2237] <= 3;
		weights[2238] <= 170;
		weights[2239] <= 192;
		weights[2240] <= 75;
		weights[2241] <= 235;
		weights[2242] <= 109;
		weights[2243] <= 27;
		weights[2244] <= 35;
		weights[2245] <= 172;
		weights[2246] <= 189;
		weights[2247] <= 15;
		weights[2248] <= 116;
		weights[2249] <= 190;
		weights[2250] <= 2;
		weights[2251] <= 49;
		weights[2252] <= 214;
		weights[2253] <= 66;
		weights[2254] <= 63;
		weights[2255] <= 1;
		weights[2256] <= 88;
		weights[2257] <= 252;
		weights[2258] <= 243;
		weights[2259] <= 61;
		weights[2260] <= 185;
		weights[2261] <= 186;
		weights[2262] <= 24;
		weights[2263] <= 219;
		weights[2264] <= 186;
		weights[2265] <= 89;
		weights[2266] <= 30;
		weights[2267] <= 187;
		weights[2268] <= 7;
		weights[2269] <= 24;
		weights[2270] <= 165;
		weights[2271] <= 101;
		weights[2272] <= 107;
		weights[2273] <= 133;
		weights[2274] <= 153;
		weights[2275] <= 12;
		weights[2276] <= 248;
		weights[2277] <= 10;
		weights[2278] <= 81;
		weights[2279] <= 106;
		weights[2280] <= 219;
		weights[2281] <= 222;
		weights[2282] <= 178;
		weights[2283] <= 86;
		weights[2284] <= 218;
		weights[2285] <= 188;
		weights[2286] <= 190;
		weights[2287] <= 232;
		weights[2288] <= 69;
		weights[2289] <= 141;
		weights[2290] <= 96;
		weights[2291] <= 244;
		weights[2292] <= 68;
		weights[2293] <= 78;
		weights[2294] <= 189;
		weights[2295] <= 212;
		weights[2296] <= 190;
		weights[2297] <= 129;
		weights[2298] <= 223;
		weights[2299] <= 138;
		weights[2300] <= 94;
		weights[2301] <= 88;
		weights[2302] <= 225;
		weights[2303] <= 157;
		weights[2304] <= 100;
		weights[2305] <= 232;
		weights[2306] <= 46;
		weights[2307] <= 20;
		weights[2308] <= 163;
		weights[2309] <= 164;
		weights[2310] <= 137;
		weights[2311] <= 55;
		weights[2312] <= 142;
		weights[2313] <= 225;
		weights[2314] <= 149;
		weights[2315] <= 97;
		weights[2316] <= 214;
		weights[2317] <= 143;
		weights[2318] <= 54;
		weights[2319] <= 74;
		weights[2320] <= 174;
		weights[2321] <= 96;
		weights[2322] <= 165;
		weights[2323] <= 81;
		weights[2324] <= 198;
		weights[2325] <= 21;
		weights[2326] <= 146;
		weights[2327] <= 4;
		weights[2328] <= 177;
		weights[2329] <= 52;
		weights[2330] <= 116;
		weights[2331] <= 156;
		weights[2332] <= 160;
		weights[2333] <= 6;
		weights[2334] <= 142;
		weights[2335] <= 95;
		weights[2336] <= 214;
		weights[2337] <= 139;
		weights[2338] <= 168;
		weights[2339] <= 39;
		weights[2340] <= 169;
		weights[2341] <= 170;
		weights[2342] <= 72;
		weights[2343] <= 106;
		weights[2344] <= 13;
		weights[2345] <= 163;
		weights[2346] <= 246;
		weights[2347] <= 113;
		weights[2348] <= 174;
		weights[2349] <= 198;
		weights[2350] <= 211;
		weights[2351] <= 121;
		weights[2352] <= 208;
		weights[2353] <= 157;
		weights[2354] <= 38;
		weights[2355] <= 164;
		weights[2356] <= 172;
		weights[2357] <= 247;
		weights[2358] <= 102;
		weights[2359] <= 51;
		weights[2360] <= 96;
		weights[2361] <= 139;
		weights[2362] <= 107;
		weights[2363] <= 200;
		weights[2364] <= 193;
		weights[2365] <= 103;
		weights[2366] <= 64;
		weights[2367] <= 117;
		weights[2368] <= 35;
		weights[2369] <= 109;
		weights[2370] <= 141;
		weights[2371] <= 35;
		weights[2372] <= 115;
		weights[2373] <= 6;
		weights[2374] <= 169;
		weights[2375] <= 83;
		weights[2376] <= 88;
		weights[2377] <= 37;
		weights[2378] <= 174;
		weights[2379] <= 33;
		weights[2380] <= 130;
		weights[2381] <= 44;
		weights[2382] <= 52;
		weights[2383] <= 103;
		weights[2384] <= 244;
		weights[2385] <= 224;
		weights[2386] <= 187;
		weights[2387] <= 50;
		weights[2388] <= 152;
		weights[2389] <= 223;
		weights[2390] <= 62;
		weights[2391] <= 222;
		weights[2392] <= 75;
		weights[2393] <= 235;
		weights[2394] <= 244;
		weights[2395] <= 75;
		weights[2396] <= 117;
		weights[2397] <= 174;
		weights[2398] <= 160;
		weights[2399] <= 23;
		weights[2400] <= 162;
		weights[2401] <= 132;
		weights[2402] <= 184;
		weights[2403] <= 49;
		weights[2404] <= 84;
		weights[2405] <= 152;
		weights[2406] <= 230;
		weights[2407] <= 249;
		weights[2408] <= 76;
		weights[2409] <= 159;
		weights[2410] <= 204;
		weights[2411] <= 117;
		weights[2412] <= 1;
		weights[2413] <= 249;
		weights[2414] <= 60;
		weights[2415] <= 221;
		weights[2416] <= 89;
		weights[2417] <= 234;
		weights[2418] <= 172;
		weights[2419] <= 166;
		weights[2420] <= 193;
		weights[2421] <= 112;
		weights[2422] <= 147;
		weights[2423] <= 61;
		weights[2424] <= 167;
		weights[2425] <= 128;
		weights[2426] <= 148;
		weights[2427] <= 141;
		weights[2428] <= 225;
		weights[2429] <= 118;
		weights[2430] <= 124;
		weights[2431] <= 75;
		weights[2432] <= 212;
		weights[2433] <= 222;
		weights[2434] <= 84;
		weights[2435] <= 238;
		weights[2436] <= 10;
		weights[2437] <= 29;
		weights[2438] <= 189;
		weights[2439] <= 158;
		weights[2440] <= 99;
		weights[2441] <= 100;
		weights[2442] <= 51;
		weights[2443] <= 251;
		weights[2444] <= 122;
		weights[2445] <= 89;
		weights[2446] <= 110;
		weights[2447] <= 246;
		weights[2448] <= 186;
		weights[2449] <= 74;
		weights[2450] <= 113;
		weights[2451] <= 227;
		weights[2452] <= 178;
		weights[2453] <= 32;
		weights[2454] <= 227;
		weights[2455] <= 228;
		weights[2456] <= 138;
		weights[2457] <= 233;
		weights[2458] <= 91;
		weights[2459] <= 210;
		weights[2460] <= 176;
		weights[2461] <= 11;
		weights[2462] <= 221;
		weights[2463] <= 39;
		weights[2464] <= 233;
		weights[2465] <= 196;
		weights[2466] <= 219;
		weights[2467] <= 184;
		weights[2468] <= 119;
		weights[2469] <= 235;
		weights[2470] <= 216;
		weights[2471] <= 144;
		weights[2472] <= 126;
		weights[2473] <= 32;
		weights[2474] <= 68;
		weights[2475] <= 109;
		weights[2476] <= 31;
		weights[2477] <= 216;
		weights[2478] <= 65;
		weights[2479] <= 126;
		weights[2480] <= 186;
		weights[2481] <= 107;
		weights[2482] <= 95;
		weights[2483] <= 237;
		weights[2484] <= 249;
		weights[2485] <= 11;
		weights[2486] <= 73;
		weights[2487] <= 228;
		weights[2488] <= 225;
		weights[2489] <= 141;
		weights[2490] <= 143;
		weights[2491] <= 229;
		weights[2492] <= 148;
		weights[2493] <= 51;
		weights[2494] <= 56;
		weights[2495] <= 77;
		weights[2496] <= 229;
		weights[2497] <= 173;
		weights[2498] <= 117;
		weights[2499] <= 132;
		weights[2500] <= 132;
		weights[2501] <= 25;
		weights[2502] <= 113;
		weights[2503] <= 203;
		weights[2504] <= 134;
		weights[2505] <= 135;
		weights[2506] <= 196;
		weights[2507] <= 100;
		weights[2508] <= 21;
		weights[2509] <= 60;
		weights[2510] <= 192;
		weights[2511] <= 72;
		weights[2512] <= 169;
		weights[2513] <= 34;
		weights[2514] <= 201;
		weights[2515] <= 138;
		weights[2516] <= 154;
		weights[2517] <= 227;
		weights[2518] <= 174;
		weights[2519] <= 219;
		weights[2520] <= 218;
		weights[2521] <= 142;
		weights[2522] <= 225;
		weights[2523] <= 137;
		weights[2524] <= 215;
		weights[2525] <= 235;
		weights[2526] <= 69;
		weights[2527] <= 227;
		weights[2528] <= 52;
		weights[2529] <= 59;
		weights[2530] <= 141;
		weights[2531] <= 62;
		weights[2532] <= 243;
		weights[2533] <= 210;
		weights[2534] <= 2;
		weights[2535] <= 255;
		weights[2536] <= 33;
		weights[2537] <= 157;
		weights[2538] <= 234;
		weights[2539] <= 36;
		weights[2540] <= 185;
		weights[2541] <= 103;
		weights[2542] <= 28;
		weights[2543] <= 176;
		weights[2544] <= 145;
		weights[2545] <= 205;
		weights[2546] <= 93;
		weights[2547] <= 80;
		weights[2548] <= 114;
		weights[2549] <= 39;
		weights[2550] <= 33;
		weights[2551] <= 93;
		weights[2552] <= 22;
		weights[2553] <= 55;
		weights[2554] <= 49;
		weights[2555] <= 183;
		weights[2556] <= 44;
		weights[2557] <= 141;
		weights[2558] <= 193;
		weights[2559] <= 107;
		weights[2560] <= 153;
		weights[2561] <= 41;
		weights[2562] <= 134;
		weights[2563] <= 82;
		weights[2564] <= 175;
		weights[2565] <= 226;
		weights[2566] <= 253;
		weights[2567] <= 107;
		weights[2568] <= 100;
		weights[2569] <= 185;
		weights[2570] <= 153;
		weights[2571] <= 187;
		weights[2572] <= 137;
		weights[2573] <= 238;
		weights[2574] <= 211;
		weights[2575] <= 181;
		weights[2576] <= 88;
		weights[2577] <= 125;
		weights[2578] <= 210;
		weights[2579] <= 110;
		weights[2580] <= 129;
		weights[2581] <= 216;
		weights[2582] <= 175;
		weights[2583] <= 193;
		weights[2584] <= 149;
		weights[2585] <= 185;
		weights[2586] <= 74;
		weights[2587] <= 201;
		weights[2588] <= 159;
		weights[2589] <= 52;
		weights[2590] <= 171;
		weights[2591] <= 163;
		weights[2592] <= 193;
		weights[2593] <= 24;
		weights[2594] <= 185;
		weights[2595] <= 64;
		weights[2596] <= 148;
		weights[2597] <= 205;
		weights[2598] <= 230;
		weights[2599] <= 127;
		weights[2600] <= 112;
		weights[2601] <= 141;
		weights[2602] <= 119;
		weights[2603] <= 222;
		weights[2604] <= 52;
		weights[2605] <= 48;
		weights[2606] <= 172;
		weights[2607] <= 88;
		weights[2608] <= 162;
		weights[2609] <= 25;
		weights[2610] <= 243;
		weights[2611] <= 69;
		weights[2612] <= 219;
		weights[2613] <= 237;
		weights[2614] <= 216;
		weights[2615] <= 163;
		weights[2616] <= 81;
		weights[2617] <= 45;
		weights[2618] <= 199;
		weights[2619] <= 238;
		weights[2620] <= 179;
		weights[2621] <= 177;
		weights[2622] <= 96;
		weights[2623] <= 147;
		weights[2624] <= 144;
		weights[2625] <= 32;
		weights[2626] <= 255;
		weights[2627] <= 47;
		weights[2628] <= 102;
		weights[2629] <= 34;
		weights[2630] <= 250;
		weights[2631] <= 224;
		weights[2632] <= 114;
		weights[2633] <= 197;
		weights[2634] <= 226;
		weights[2635] <= 151;
		weights[2636] <= 48;
		weights[2637] <= 253;
		weights[2638] <= 34;
		weights[2639] <= 128;
		weights[2640] <= 20;
		weights[2641] <= 235;
		weights[2642] <= 158;
		weights[2643] <= 116;
		weights[2644] <= 113;
		weights[2645] <= 86;
		weights[2646] <= 239;
		weights[2647] <= 235;
		weights[2648] <= 103;
		weights[2649] <= 208;
		weights[2650] <= 197;
		weights[2651] <= 137;
		weights[2652] <= 120;
		weights[2653] <= 251;
		weights[2654] <= 16;
		weights[2655] <= 55;
		weights[2656] <= 48;
		weights[2657] <= 163;
		weights[2658] <= 5;
		weights[2659] <= 94;
		weights[2660] <= 131;
		weights[2661] <= 178;
		weights[2662] <= 170;
		weights[2663] <= 230;
		weights[2664] <= 82;
		weights[2665] <= 35;
		weights[2666] <= 207;
		weights[2667] <= 193;
		weights[2668] <= 224;
		weights[2669] <= 77;
		weights[2670] <= 124;
		weights[2671] <= 34;
		weights[2672] <= 82;
		weights[2673] <= 216;
		weights[2674] <= 37;
		weights[2675] <= 203;
		weights[2676] <= 105;
		weights[2677] <= 218;
		weights[2678] <= 74;
		weights[2679] <= 181;
		weights[2680] <= 52;
		weights[2681] <= 243;
		weights[2682] <= 165;
		weights[2683] <= 45;
		weights[2684] <= 50;
		weights[2685] <= 199;
		weights[2686] <= 19;
		weights[2687] <= 204;
		weights[2688] <= 110;
		weights[2689] <= 11;
		weights[2690] <= 12;
		weights[2691] <= 176;
		weights[2692] <= 88;
		weights[2693] <= 167;
		weights[2694] <= 48;
		weights[2695] <= 152;
		weights[2696] <= 189;
		weights[2697] <= 77;
		weights[2698] <= 125;
		weights[2699] <= 193;
		weights[2700] <= 181;
		weights[2701] <= 107;
		weights[2702] <= 240;
		weights[2703] <= 36;
		weights[2704] <= 234;
		weights[2705] <= 21;
		weights[2706] <= 243;
		weights[2707] <= 64;
		weights[2708] <= 239;
		weights[2709] <= 147;
		weights[2710] <= 44;
		weights[2711] <= 250;
		weights[2712] <= 214;
		weights[2713] <= 171;
		weights[2714] <= 175;
		weights[2715] <= 135;
		weights[2716] <= 110;
		weights[2717] <= 173;
		weights[2718] <= 216;
		weights[2719] <= 241;
		weights[2720] <= 23;
		weights[2721] <= 188;
		weights[2722] <= 148;
		weights[2723] <= 78;
		weights[2724] <= 144;
		weights[2725] <= 227;
		weights[2726] <= 166;
		weights[2727] <= 154;
		weights[2728] <= 121;
		weights[2729] <= 160;
		weights[2730] <= 192;
		weights[2731] <= 190;
		weights[2732] <= 234;
		weights[2733] <= 239;
		weights[2734] <= 15;
		weights[2735] <= 57;
		weights[2736] <= 129;
		weights[2737] <= 118;
		weights[2738] <= 125;
		weights[2739] <= 16;
		weights[2740] <= 234;
		weights[2741] <= 115;
		weights[2742] <= 33;
		weights[2743] <= 46;
		weights[2744] <= 174;
		weights[2745] <= 37;
		weights[2746] <= 20;
		weights[2747] <= 156;
		weights[2748] <= 248;
		weights[2749] <= 194;
		weights[2750] <= 43;
		weights[2751] <= 46;
		weights[2752] <= 115;
		weights[2753] <= 211;
		weights[2754] <= 239;
		weights[2755] <= 44;
		weights[2756] <= 30;
		weights[2757] <= 95;
		weights[2758] <= 88;
		weights[2759] <= 161;
		weights[2760] <= 41;
		weights[2761] <= 141;
		weights[2762] <= 18;
		weights[2763] <= 175;
		weights[2764] <= 23;
		weights[2765] <= 183;
		weights[2766] <= 47;
		weights[2767] <= 39;
		weights[2768] <= 73;
		weights[2769] <= 33;
		weights[2770] <= 161;
		weights[2771] <= 56;
		weights[2772] <= 193;
		weights[2773] <= 68;
		weights[2774] <= 204;
		weights[2775] <= 14;
		weights[2776] <= 102;
		weights[2777] <= 43;
		weights[2778] <= 91;
		weights[2779] <= 136;
		weights[2780] <= 116;
		weights[2781] <= 195;
		weights[2782] <= 195;
		weights[2783] <= 86;
		weights[2784] <= 162;
		weights[2785] <= 125;
		weights[2786] <= 254;
		weights[2787] <= 98;
		weights[2788] <= 234;
		weights[2789] <= 225;
		weights[2790] <= 134;
		weights[2791] <= 140;
		weights[2792] <= 65;
		weights[2793] <= 150;
		weights[2794] <= 71;
		weights[2795] <= 121;
		weights[2796] <= 197;
		weights[2797] <= 2;
		weights[2798] <= 102;
		weights[2799] <= 225;
		weights[2800] <= 233;
		weights[2801] <= 54;
		weights[2802] <= 93;
		weights[2803] <= 78;
		weights[2804] <= 75;
		weights[2805] <= 74;
		weights[2806] <= 110;
		weights[2807] <= 93;
		weights[2808] <= 184;
		weights[2809] <= 79;
		weights[2810] <= 226;
		weights[2811] <= 125;
		weights[2812] <= 240;
		weights[2813] <= 189;
		weights[2814] <= 220;
		weights[2815] <= 243;
		weights[2816] <= 163;
		weights[2817] <= 188;
		weights[2818] <= 222;
		weights[2819] <= 126;
		weights[2820] <= 144;
		weights[2821] <= 196;
		weights[2822] <= 84;
		weights[2823] <= 90;
		weights[2824] <= 212;
		weights[2825] <= 4;
		weights[2826] <= 4;
		weights[2827] <= 90;
		weights[2828] <= 172;
		weights[2829] <= 106;
		weights[2830] <= 206;
		weights[2831] <= 248;
		weights[2832] <= 24;
		weights[2833] <= 238;
		weights[2834] <= 76;
		weights[2835] <= 56;
		weights[2836] <= 115;
		weights[2837] <= 199;
		weights[2838] <= 67;
		weights[2839] <= 245;
		weights[2840] <= 26;
		weights[2841] <= 14;
		weights[2842] <= 8;
		weights[2843] <= 135;
		weights[2844] <= 29;
		weights[2845] <= 234;
		weights[2846] <= 113;
		weights[2847] <= 41;
		weights[2848] <= 95;
		weights[2849] <= 228;
		weights[2850] <= 212;
		weights[2851] <= 197;
		weights[2852] <= 244;
		weights[2853] <= 131;
		weights[2854] <= 30;
		weights[2855] <= 196;
		weights[2856] <= 8;
		weights[2857] <= 198;
		weights[2858] <= 224;
		weights[2859] <= 177;
		weights[2860] <= 167;
		weights[2861] <= 197;
		weights[2862] <= 219;
		weights[2863] <= 158;
		weights[2864] <= 174;
		weights[2865] <= 174;
		weights[2866] <= 251;
		weights[2867] <= 218;
		weights[2868] <= 131;
		weights[2869] <= 37;
		weights[2870] <= 126;
		weights[2871] <= 104;
		weights[2872] <= 199;
		weights[2873] <= 38;
		weights[2874] <= 240;
		weights[2875] <= 197;
		weights[2876] <= 50;
		weights[2877] <= 160;
		weights[2878] <= 109;
		weights[2879] <= 183;
		weights[2880] <= 188;
		weights[2881] <= 65;
		weights[2882] <= 224;
		weights[2883] <= 122;
		weights[2884] <= 85;
		weights[2885] <= 25;
		weights[2886] <= 142;
		weights[2887] <= 86;
		weights[2888] <= 159;
		weights[2889] <= 151;
		weights[2890] <= 106;
		weights[2891] <= 115;
		weights[2892] <= 33;
		weights[2893] <= 203;
		weights[2894] <= 58;
		weights[2895] <= 24;
		weights[2896] <= 112;
		weights[2897] <= 19;
		weights[2898] <= 140;
		weights[2899] <= 67;
		weights[2900] <= 241;
		weights[2901] <= 212;
		weights[2902] <= 122;
		weights[2903] <= 12;
		weights[2904] <= 128;
		weights[2905] <= 83;
		weights[2906] <= 112;
		weights[2907] <= 140;
		weights[2908] <= 216;
		weights[2909] <= 54;
		weights[2910] <= 136;
		weights[2911] <= 23;
		weights[2912] <= 254;
		weights[2913] <= 152;
		weights[2914] <= 254;
		weights[2915] <= 118;
		weights[2916] <= 216;
		weights[2917] <= 159;
		weights[2918] <= 240;
		weights[2919] <= 111;
		weights[2920] <= 50;
		weights[2921] <= 232;
		weights[2922] <= 231;
		weights[2923] <= 95;
		weights[2924] <= 33;
		weights[2925] <= 15;
		weights[2926] <= 198;
		weights[2927] <= 58;
		weights[2928] <= 16;
		weights[2929] <= 222;
		weights[2930] <= 88;
		weights[2931] <= 194;
		weights[2932] <= 46;
		weights[2933] <= 150;
		weights[2934] <= 107;
		weights[2935] <= 120;
		weights[2936] <= 182;
		weights[2937] <= 28;
		weights[2938] <= 139;
		weights[2939] <= 26;
		weights[2940] <= 216;
		weights[2941] <= 97;
		weights[2942] <= 36;
		weights[2943] <= 128;
		weights[2944] <= 106;
		weights[2945] <= 245;
		weights[2946] <= 167;
		weights[2947] <= 68;
		weights[2948] <= 158;
		weights[2949] <= 12;
		weights[2950] <= 136;
		weights[2951] <= 185;
		weights[2952] <= 218;
		weights[2953] <= 80;
		weights[2954] <= 220;
		weights[2955] <= 58;
		weights[2956] <= 150;
		weights[2957] <= 10;
		weights[2958] <= 72;
		weights[2959] <= 113;
		weights[2960] <= 92;
		weights[2961] <= 19;
		weights[2962] <= 68;
		weights[2963] <= 26;
		weights[2964] <= 95;
		weights[2965] <= 8;
		weights[2966] <= 78;
		weights[2967] <= 226;
		weights[2968] <= 13;
		weights[2969] <= 161;
		weights[2970] <= 118;
		weights[2971] <= 65;
		weights[2972] <= 226;
		weights[2973] <= 103;
		weights[2974] <= 212;
		weights[2975] <= 93;
		weights[2976] <= 244;
		weights[2977] <= 35;
		weights[2978] <= 228;
		weights[2979] <= 237;
		weights[2980] <= 193;
		weights[2981] <= 63;
		weights[2982] <= 96;
		weights[2983] <= 89;
		weights[2984] <= 121;
		weights[2985] <= 223;
		weights[2986] <= 16;
		weights[2987] <= 102;
		weights[2988] <= 35;
		weights[2989] <= 192;
		weights[2990] <= 158;
		weights[2991] <= 226;
		weights[2992] <= 131;
		weights[2993] <= 140;
		weights[2994] <= 71;
		weights[2995] <= 166;
		weights[2996] <= 92;
		weights[2997] <= 192;
		weights[2998] <= 122;
		weights[2999] <= 161;
		weights[3000] <= 10;
		weights[3001] <= 217;
		weights[3002] <= 72;
		weights[3003] <= 221;
		weights[3004] <= 216;
		weights[3005] <= 210;
		weights[3006] <= 51;
		weights[3007] <= 209;
		weights[3008] <= 42;
		weights[3009] <= 75;
		weights[3010] <= 114;
		weights[3011] <= 35;
		weights[3012] <= 191;
		weights[3013] <= 193;
		weights[3014] <= 118;
		weights[3015] <= 253;
		weights[3016] <= 52;
		weights[3017] <= 92;
		weights[3018] <= 189;
		weights[3019] <= 220;
		weights[3020] <= 33;
		weights[3021] <= 223;
		weights[3022] <= 85;
		weights[3023] <= 9;
		weights[3024] <= 93;
		weights[3025] <= 130;
		weights[3026] <= 144;
		weights[3027] <= 218;
		weights[3028] <= 242;
		weights[3029] <= 212;
		weights[3030] <= 186;
		weights[3031] <= 224;
		weights[3032] <= 125;
		weights[3033] <= 139;
		weights[3034] <= 15;
		weights[3035] <= 21;
		weights[3036] <= 68;
		weights[3037] <= 43;
		weights[3038] <= 90;
		weights[3039] <= 230;
		weights[3040] <= 84;
		weights[3041] <= 157;
		weights[3042] <= 254;
		weights[3043] <= 154;
		weights[3044] <= 50;
		weights[3045] <= 123;
		weights[3046] <= 14;
		weights[3047] <= 185;
		weights[3048] <= 151;
		weights[3049] <= 64;
		weights[3050] <= 182;
		weights[3051] <= 11;
		weights[3052] <= 45;
		weights[3053] <= 103;
		weights[3054] <= 33;
		weights[3055] <= 91;
		weights[3056] <= 22;
		weights[3057] <= 173;
		weights[3058] <= 167;
		weights[3059] <= 33;
		weights[3060] <= 54;
		weights[3061] <= 243;
		weights[3062] <= 17;
		weights[3063] <= 151;
		weights[3064] <= 115;
		weights[3065] <= 240;
		weights[3066] <= 83;
		weights[3067] <= 224;
		weights[3068] <= 220;
		weights[3069] <= 163;
		weights[3070] <= 73;
		weights[3071] <= 121;
		weights[3072] <= 114;
		weights[3073] <= 215;
		weights[3074] <= 111;
		weights[3075] <= 143;
		weights[3076] <= 132;
		weights[3077] <= 26;
		weights[3078] <= 82;
		weights[3079] <= 192;
		weights[3080] <= 63;
		weights[3081] <= 87;
		weights[3082] <= 25;
		weights[3083] <= 151;
		weights[3084] <= 229;
		weights[3085] <= 135;
		weights[3086] <= 48;
		weights[3087] <= 47;
		weights[3088] <= 5;
		weights[3089] <= 103;
		weights[3090] <= 200;
		weights[3091] <= 38;
		weights[3092] <= 138;
		weights[3093] <= 18;
		weights[3094] <= 158;
		weights[3095] <= 35;
		weights[3096] <= 151;
		weights[3097] <= 55;
		weights[3098] <= 149;
		weights[3099] <= 16;
		weights[3100] <= 221;
		weights[3101] <= 181;
		weights[3102] <= 31;
		weights[3103] <= 27;
		weights[3104] <= 172;
		weights[3105] <= 235;
		weights[3106] <= 228;
		weights[3107] <= 232;
		weights[3108] <= 182;
		weights[3109] <= 218;
		weights[3110] <= 149;
		weights[3111] <= 39;
		weights[3112] <= 210;
		weights[3113] <= 214;
		weights[3114] <= 242;
		weights[3115] <= 211;
		weights[3116] <= 133;
		weights[3117] <= 115;
		weights[3118] <= 82;
		weights[3119] <= 72;
		weights[3120] <= 170;
		weights[3121] <= 44;
		weights[3122] <= 219;
		weights[3123] <= 99;
		weights[3124] <= 145;
		weights[3125] <= 148;
		weights[3126] <= 50;
		weights[3127] <= 133;
		weights[3128] <= 241;
		weights[3129] <= 145;
		weights[3130] <= 1;
		weights[3131] <= 178;
		weights[3132] <= 191;
		weights[3133] <= 110;
		weights[3134] <= 238;
		weights[3135] <= 101;
		weights[3136] <= 29;
		weights[3137] <= 17;
		weights[3138] <= 39;
		weights[3139] <= 68;
		weights[3140] <= 68;
		weights[3141] <= 234;
		weights[3142] <= 103;
		weights[3143] <= 222;
		weights[3144] <= 73;
		weights[3145] <= 219;
		weights[3146] <= 228;
		weights[3147] <= 237;
		weights[3148] <= 87;
		weights[3149] <= 13;
		weights[3150] <= 44;
		weights[3151] <= 249;
		weights[3152] <= 115;
		weights[3153] <= 219;
		weights[3154] <= 204;
		weights[3155] <= 250;
		weights[3156] <= 22;
		weights[3157] <= 145;
		weights[3158] <= 75;
		weights[3159] <= 94;
		weights[3160] <= 82;
		weights[3161] <= 70;
		weights[3162] <= 62;
		weights[3163] <= 246;
		weights[3164] <= 49;
		weights[3165] <= 186;
		weights[3166] <= 108;
		weights[3167] <= 69;
		weights[3168] <= 155;
		weights[3169] <= 13;
		weights[3170] <= 249;
		weights[3171] <= 18;
		weights[3172] <= 161;
		weights[3173] <= 91;
		weights[3174] <= 36;
		weights[3175] <= 161;
		weights[3176] <= 241;
		weights[3177] <= 38;
		weights[3178] <= 140;
		weights[3179] <= 134;
		weights[3180] <= 183;
		weights[3181] <= 32;
		weights[3182] <= 128;
		weights[3183] <= 54;
		weights[3184] <= 50;
		weights[3185] <= 123;
		weights[3186] <= 121;
		weights[3187] <= 100;
		weights[3188] <= 54;
		weights[3189] <= 82;
		weights[3190] <= 235;
		weights[3191] <= 170;
		weights[3192] <= 241;
		weights[3193] <= 104;
		weights[3194] <= 207;
		weights[3195] <= 146;
		weights[3196] <= 211;
		weights[3197] <= 2;
		weights[3198] <= 129;
		weights[3199] <= 184;
		weights[3200] <= 233;
		weights[3201] <= 107;
		weights[3202] <= 123;
		weights[3203] <= 203;
		weights[3204] <= 89;
		weights[3205] <= 14;
		weights[3206] <= 191;
		weights[3207] <= 55;
		weights[3208] <= 62;
		weights[3209] <= 172;
		weights[3210] <= 227;
		weights[3211] <= 3;
		weights[3212] <= 122;
		weights[3213] <= 178;
		weights[3214] <= 91;
		weights[3215] <= 67;
		weights[3216] <= 55;
		weights[3217] <= 184;
		weights[3218] <= 218;
		weights[3219] <= 176;
		weights[3220] <= 233;
		weights[3221] <= 203;
		weights[3222] <= 236;
		weights[3223] <= 224;
		weights[3224] <= 84;
		weights[3225] <= 122;
		weights[3226] <= 14;
		weights[3227] <= 205;
		weights[3228] <= 23;
		weights[3229] <= 78;
		weights[3230] <= 29;
		weights[3231] <= 207;
		weights[3232] <= 238;
		weights[3233] <= 100;
		weights[3234] <= 61;
		weights[3235] <= 61;
		weights[3236] <= 47;
		weights[3237] <= 218;
		weights[3238] <= 82;
		weights[3239] <= 186;
		weights[3240] <= 43;
		weights[3241] <= 36;
		weights[3242] <= 208;
		weights[3243] <= 194;
		weights[3244] <= 173;
		weights[3245] <= 183;
		weights[3246] <= 166;
		weights[3247] <= 164;
		weights[3248] <= 203;
		weights[3249] <= 206;
		weights[3250] <= 79;
		weights[3251] <= 155;
		weights[3252] <= 238;
		weights[3253] <= 20;
		weights[3254] <= 201;
		weights[3255] <= 108;
		weights[3256] <= 152;
		weights[3257] <= 130;
		weights[3258] <= 13;
		weights[3259] <= 228;
		weights[3260] <= 75;
		weights[3261] <= 46;
		weights[3262] <= 93;
		weights[3263] <= 203;
		weights[3264] <= 235;
		weights[3265] <= 100;
		weights[3266] <= 238;
		weights[3267] <= 22;
		weights[3268] <= 121;
		weights[3269] <= 229;
		weights[3270] <= 99;
		weights[3271] <= 220;
		weights[3272] <= 253;
		weights[3273] <= 206;
		weights[3274] <= 70;
		weights[3275] <= 209;
		weights[3276] <= 51;
		weights[3277] <= 117;
		weights[3278] <= 73;
		weights[3279] <= 108;
		weights[3280] <= 72;
		weights[3281] <= 196;
		weights[3282] <= 100;
		weights[3283] <= 39;
		weights[3284] <= 102;
		weights[3285] <= 160;
		weights[3286] <= 232;
		weights[3287] <= 40;
		weights[3288] <= 124;
		weights[3289] <= 218;
		weights[3290] <= 85;
		weights[3291] <= 69;
		weights[3292] <= 130;
		weights[3293] <= 115;
		weights[3294] <= 89;
		weights[3295] <= 5;
		weights[3296] <= 13;
		weights[3297] <= 155;
		weights[3298] <= 88;
		weights[3299] <= 185;
		weights[3300] <= 82;
		weights[3301] <= 28;
		weights[3302] <= 16;
		weights[3303] <= 246;
		weights[3304] <= 161;
		weights[3305] <= 61;
		weights[3306] <= 96;
		weights[3307] <= 249;
		weights[3308] <= 42;
		weights[3309] <= 68;
		weights[3310] <= 108;
		weights[3311] <= 200;
		weights[3312] <= 112;
		weights[3313] <= 57;
		weights[3314] <= 184;
		weights[3315] <= 224;
		weights[3316] <= 80;
		weights[3317] <= 235;
		weights[3318] <= 50;
		weights[3319] <= 219;
		weights[3320] <= 238;
		weights[3321] <= 253;
		weights[3322] <= 169;
		weights[3323] <= 201;
		weights[3324] <= 26;
		weights[3325] <= 82;
		weights[3326] <= 237;
		weights[3327] <= 119;
		weights[3328] <= 71;
		weights[3329] <= 244;
		weights[3330] <= 102;
		weights[3331] <= 35;
		weights[3332] <= 249;
		weights[3333] <= 40;
		weights[3334] <= 95;
		weights[3335] <= 6;
		weights[3336] <= 252;
		weights[3337] <= 128;
		weights[3338] <= 20;
		weights[3339] <= 12;
		weights[3340] <= 5;
		weights[3341] <= 127;
		weights[3342] <= 10;
		weights[3343] <= 143;
		weights[3344] <= 70;
		weights[3345] <= 214;
		weights[3346] <= 233;
		weights[3347] <= 103;
		weights[3348] <= 126;
		weights[3349] <= 241;
		weights[3350] <= 244;
		weights[3351] <= 76;
		weights[3352] <= 76;
		weights[3353] <= 114;
		weights[3354] <= 5;
		weights[3355] <= 49;
		weights[3356] <= 32;
		weights[3357] <= 185;
		weights[3358] <= 67;
		weights[3359] <= 83;
		weights[3360] <= 106;
		weights[3361] <= 45;
		weights[3362] <= 19;
		weights[3363] <= 115;
		weights[3364] <= 134;
		weights[3365] <= 167;
		weights[3366] <= 218;
		weights[3367] <= 141;
		weights[3368] <= 224;
		weights[3369] <= 96;
		weights[3370] <= 57;
		weights[3371] <= 68;
		weights[3372] <= 232;
		weights[3373] <= 121;
		weights[3374] <= 255;
		weights[3375] <= 156;
		weights[3376] <= 9;
		weights[3377] <= 79;
		weights[3378] <= 32;
		weights[3379] <= 216;
		weights[3380] <= 55;
		weights[3381] <= 118;
		weights[3382] <= 115;
		weights[3383] <= 13;
		weights[3384] <= 235;
		weights[3385] <= 221;
		weights[3386] <= 200;
		weights[3387] <= 54;
		weights[3388] <= 206;
		weights[3389] <= 89;
		weights[3390] <= 220;
		weights[3391] <= 154;
		weights[3392] <= 98;
		weights[3393] <= 179;
		weights[3394] <= 220;
		weights[3395] <= 44;
		weights[3396] <= 140;
		weights[3397] <= 164;
		weights[3398] <= 211;
		weights[3399] <= 129;
		weights[3400] <= 55;
		weights[3401] <= 208;
		weights[3402] <= 108;
		weights[3403] <= 248;
		weights[3404] <= 17;
		weights[3405] <= 232;
		weights[3406] <= 157;
		weights[3407] <= 115;
		weights[3408] <= 227;
		weights[3409] <= 216;
		weights[3410] <= 139;
		weights[3411] <= 40;
		weights[3412] <= 57;
		weights[3413] <= 21;
		weights[3414] <= 154;
		weights[3415] <= 59;
		weights[3416] <= 29;
		weights[3417] <= 134;
		weights[3418] <= 100;
		weights[3419] <= 225;
		weights[3420] <= 215;
		weights[3421] <= 92;
		weights[3422] <= 106;
		weights[3423] <= 126;
		weights[3424] <= 36;
		weights[3425] <= 223;
		weights[3426] <= 218;
		weights[3427] <= 183;
		weights[3428] <= 38;
		weights[3429] <= 89;
		weights[3430] <= 194;
		weights[3431] <= 51;
		weights[3432] <= 197;
		weights[3433] <= 109;
		weights[3434] <= 144;
		weights[3435] <= 163;
		weights[3436] <= 115;
		weights[3437] <= 170;
		weights[3438] <= 65;
		weights[3439] <= 93;
		weights[3440] <= 215;
		weights[3441] <= 27;
		weights[3442] <= 235;
		weights[3443] <= 165;
		weights[3444] <= 239;
		weights[3445] <= 24;
		weights[3446] <= 116;
		weights[3447] <= 252;
		weights[3448] <= 94;
		weights[3449] <= 186;
		weights[3450] <= 182;
		weights[3451] <= 241;
		weights[3452] <= 223;
		weights[3453] <= 50;
		weights[3454] <= 142;
		weights[3455] <= 101;
		weights[3456] <= 216;
		weights[3457] <= 171;
		weights[3458] <= 211;
		weights[3459] <= 129;
		weights[3460] <= 171;
		weights[3461] <= 242;
		weights[3462] <= 206;
		weights[3463] <= 237;
		weights[3464] <= 203;
		weights[3465] <= 117;
		weights[3466] <= 27;
		weights[3467] <= 95;
		weights[3468] <= 192;
		weights[3469] <= 232;
		weights[3470] <= 79;
		weights[3471] <= 184;
		weights[3472] <= 252;
		weights[3473] <= 174;
		weights[3474] <= 160;
		weights[3475] <= 43;
		weights[3476] <= 173;
		weights[3477] <= 178;
		weights[3478] <= 140;
		weights[3479] <= 177;
		weights[3480] <= 186;
		weights[3481] <= 94;
		weights[3482] <= 6;
		weights[3483] <= 19;
		weights[3484] <= 77;
		weights[3485] <= 181;
		weights[3486] <= 168;
		weights[3487] <= 131;
		weights[3488] <= 188;
		weights[3489] <= 141;
		weights[3490] <= 199;
		weights[3491] <= 204;
		weights[3492] <= 207;
		weights[3493] <= 193;
		weights[3494] <= 178;
		weights[3495] <= 138;
		weights[3496] <= 34;
		weights[3497] <= 40;
		weights[3498] <= 100;
		weights[3499] <= 49;
		weights[3500] <= 152;
		weights[3501] <= 33;
		weights[3502] <= 237;
		weights[3503] <= 146;
		weights[3504] <= 101;
		weights[3505] <= 247;
		weights[3506] <= 203;
		weights[3507] <= 172;
		weights[3508] <= 161;
		weights[3509] <= 51;
		weights[3510] <= 196;
		weights[3511] <= 50;
		weights[3512] <= 197;
		weights[3513] <= 230;
		weights[3514] <= 195;
		weights[3515] <= 219;
		weights[3516] <= 212;
		weights[3517] <= 196;
		weights[3518] <= 6;
		weights[3519] <= 119;
		weights[3520] <= 144;
		weights[3521] <= 44;
		weights[3522] <= 253;
		weights[3523] <= 93;
		weights[3524] <= 204;
		weights[3525] <= 54;
		weights[3526] <= 26;
		weights[3527] <= 8;
		weights[3528] <= 78;
		weights[3529] <= 36;
		weights[3530] <= 194;
		weights[3531] <= 8;
		weights[3532] <= 95;
		weights[3533] <= 193;
		weights[3534] <= 194;
		weights[3535] <= 57;
		weights[3536] <= 232;
		weights[3537] <= 54;
		weights[3538] <= 5;
		weights[3539] <= 157;
		weights[3540] <= 111;
		weights[3541] <= 200;
		weights[3542] <= 168;
		weights[3543] <= 214;
		weights[3544] <= 171;
		weights[3545] <= 48;
		weights[3546] <= 8;
		weights[3547] <= 95;
		weights[3548] <= 105;
		weights[3549] <= 85;
		weights[3550] <= 53;
		weights[3551] <= 129;
		weights[3552] <= 35;
		weights[3553] <= 20;
		weights[3554] <= 185;
		weights[3555] <= 90;
		weights[3556] <= 7;
		weights[3557] <= 225;
		weights[3558] <= 22;
		weights[3559] <= 87;
		weights[3560] <= 18;
		weights[3561] <= 86;
		weights[3562] <= 116;
		weights[3563] <= 131;
		weights[3564] <= 147;
		weights[3565] <= 129;
		weights[3566] <= 214;
		weights[3567] <= 215;
		weights[3568] <= 104;
		weights[3569] <= 164;
		weights[3570] <= 180;
		weights[3571] <= 63;
		weights[3572] <= 250;
		weights[3573] <= 165;
		weights[3574] <= 29;
		weights[3575] <= 150;
		weights[3576] <= 80;
		weights[3577] <= 213;
		weights[3578] <= 23;
		weights[3579] <= 172;
		weights[3580] <= 37;
		weights[3581] <= 3;
		weights[3582] <= 73;
		weights[3583] <= 89;
		weights[3584] <= 81;
		weights[3585] <= 241;
		weights[3586] <= 205;
		weights[3587] <= 94;
		weights[3588] <= 10;
		weights[3589] <= 156;
		weights[3590] <= 166;
		weights[3591] <= 195;
		weights[3592] <= 221;
		weights[3593] <= 151;
		weights[3594] <= 117;
		weights[3595] <= 75;
		weights[3596] <= 131;
		weights[3597] <= 126;
		weights[3598] <= 116;
		weights[3599] <= 140;
		weights[3600] <= 50;
		weights[3601] <= 111;
		weights[3602] <= 206;
		weights[3603] <= 95;
		weights[3604] <= 157;
		weights[3605] <= 233;
		weights[3606] <= 10;
		weights[3607] <= 216;
		weights[3608] <= 112;
		weights[3609] <= 116;
		weights[3610] <= 106;
		weights[3611] <= 99;
		weights[3612] <= 217;
		weights[3613] <= 132;
		weights[3614] <= 167;
		weights[3615] <= 211;
		weights[3616] <= 133;
		weights[3617] <= 163;
		weights[3618] <= 80;
		weights[3619] <= 120;
		weights[3620] <= 1;
		weights[3621] <= 148;
		weights[3622] <= 112;
		weights[3623] <= 111;
		weights[3624] <= 131;
		weights[3625] <= 92;
		weights[3626] <= 41;
		weights[3627] <= 12;
		weights[3628] <= 223;
		weights[3629] <= 114;
		weights[3630] <= 191;
		weights[3631] <= 135;
		weights[3632] <= 184;
		weights[3633] <= 218;
		weights[3634] <= 65;
		weights[3635] <= 61;
		weights[3636] <= 190;
		weights[3637] <= 103;
		weights[3638] <= 223;
		weights[3639] <= 202;
		weights[3640] <= 13;
		weights[3641] <= 76;
		weights[3642] <= 55;
		weights[3643] <= 96;
		weights[3644] <= 23;
		weights[3645] <= 146;
		weights[3646] <= 96;
		weights[3647] <= 174;
		weights[3648] <= 27;
		weights[3649] <= 168;
		weights[3650] <= 37;
		weights[3651] <= 82;
		weights[3652] <= 225;
		weights[3653] <= 115;
		weights[3654] <= 61;
		weights[3655] <= 76;
		weights[3656] <= 152;
		weights[3657] <= 240;
		weights[3658] <= 247;
		weights[3659] <= 30;
		weights[3660] <= 174;
		weights[3661] <= 194;
		weights[3662] <= 215;
		weights[3663] <= 12;
		weights[3664] <= 94;
		weights[3665] <= 163;
		weights[3666] <= 88;
		weights[3667] <= 60;
		weights[3668] <= 157;
		weights[3669] <= 78;
		weights[3670] <= 32;
		weights[3671] <= 190;
		weights[3672] <= 242;
		weights[3673] <= 29;
		weights[3674] <= 33;
		weights[3675] <= 226;
		weights[3676] <= 14;
		weights[3677] <= 24;
		weights[3678] <= 140;
		weights[3679] <= 178;
		weights[3680] <= 248;
		weights[3681] <= 199;
		weights[3682] <= 224;
		weights[3683] <= 71;
		weights[3684] <= 174;
		weights[3685] <= 145;
		weights[3686] <= 58;
		weights[3687] <= 138;
		weights[3688] <= 12;
		weights[3689] <= 56;
		weights[3690] <= 181;
		weights[3691] <= 190;
		weights[3692] <= 169;
		weights[3693] <= 78;
		weights[3694] <= 27;
		weights[3695] <= 93;
		weights[3696] <= 35;
		weights[3697] <= 173;
		weights[3698] <= 177;
		weights[3699] <= 142;
		weights[3700] <= 31;
		weights[3701] <= 240;
		weights[3702] <= 235;
		weights[3703] <= 221;
		weights[3704] <= 129;
		weights[3705] <= 105;
		weights[3706] <= 210;
		weights[3707] <= 168;
		weights[3708] <= 220;
		weights[3709] <= 123;
		weights[3710] <= 233;
		weights[3711] <= 156;
		weights[3712] <= 90;
		weights[3713] <= 109;
		weights[3714] <= 45;
		weights[3715] <= 101;
		weights[3716] <= 124;
		weights[3717] <= 56;
		weights[3718] <= 255;
		weights[3719] <= 85;
		weights[3720] <= 59;
		weights[3721] <= 23;
		weights[3722] <= 228;
		weights[3723] <= 208;
		weights[3724] <= 148;
		weights[3725] <= 203;
		weights[3726] <= 44;
		weights[3727] <= 178;
		weights[3728] <= 130;
		weights[3729] <= 254;
		weights[3730] <= 163;
		weights[3731] <= 32;
		weights[3732] <= 42;
		weights[3733] <= 105;
		weights[3734] <= 224;
		weights[3735] <= 193;
		weights[3736] <= 3;
		weights[3737] <= 243;
		weights[3738] <= 42;
		weights[3739] <= 32;
		weights[3740] <= 216;
		weights[3741] <= 225;
		weights[3742] <= 182;
		weights[3743] <= 56;
		weights[3744] <= 160;
		weights[3745] <= 128;
		weights[3746] <= 59;
		weights[3747] <= 224;
		weights[3748] <= 25;
		weights[3749] <= 204;
		weights[3750] <= 111;
		weights[3751] <= 45;
		weights[3752] <= 63;
		weights[3753] <= 183;
		weights[3754] <= 36;
		weights[3755] <= 167;
		weights[3756] <= 84;
		weights[3757] <= 200;
		weights[3758] <= 154;
		weights[3759] <= 72;
		weights[3760] <= 208;
		weights[3761] <= 69;
		weights[3762] <= 172;
		weights[3763] <= 189;
		weights[3764] <= 135;
		weights[3765] <= 208;
		weights[3766] <= 209;
		weights[3767] <= 166;
		weights[3768] <= 205;
		weights[3769] <= 161;
		weights[3770] <= 166;
		weights[3771] <= 54;
		weights[3772] <= 221;
		weights[3773] <= 219;
		weights[3774] <= 75;
		weights[3775] <= 117;
		weights[3776] <= 241;
		weights[3777] <= 149;
		weights[3778] <= 50;
		weights[3779] <= 237;
		weights[3780] <= 73;
		weights[3781] <= 4;
		weights[3782] <= 250;
		weights[3783] <= 236;
		weights[3784] <= 102;
		weights[3785] <= 6;
		weights[3786] <= 142;
		weights[3787] <= 133;
		weights[3788] <= 127;
		weights[3789] <= 167;
		weights[3790] <= 108;
		weights[3791] <= 188;
		weights[3792] <= 156;
		weights[3793] <= 241;
		weights[3794] <= 33;
		weights[3795] <= 231;
		weights[3796] <= 145;
		weights[3797] <= 16;
		weights[3798] <= 113;
		weights[3799] <= 129;
		weights[3800] <= 65;
		weights[3801] <= 100;
		weights[3802] <= 203;
		weights[3803] <= 108;
		weights[3804] <= 181;
		weights[3805] <= 151;
		weights[3806] <= 18;
		weights[3807] <= 69;
		weights[3808] <= 200;
		weights[3809] <= 93;
		weights[3810] <= 160;
		weights[3811] <= 110;
		weights[3812] <= 102;
		weights[3813] <= 229;
		weights[3814] <= 16;
		weights[3815] <= 238;
		weights[3816] <= 41;
		weights[3817] <= 94;
		weights[3818] <= 209;
		weights[3819] <= 193;
		weights[3820] <= 14;
		weights[3821] <= 186;
		weights[3822] <= 67;
		weights[3823] <= 34;
		weights[3824] <= 103;
		weights[3825] <= 200;
		weights[3826] <= 228;
		weights[3827] <= 103;
		weights[3828] <= 227;
		weights[3829] <= 255;
		weights[3830] <= 74;
		weights[3831] <= 29;
		weights[3832] <= 150;
		weights[3833] <= 169;
		weights[3834] <= 11;
		weights[3835] <= 59;
		weights[3836] <= 52;
		weights[3837] <= 7;
		weights[3838] <= 103;
		weights[3839] <= 101;
		weights[3840] <= 177;
		weights[3841] <= 19;
		weights[3842] <= 35;
		weights[3843] <= 57;
		weights[3844] <= 248;
		weights[3845] <= 16;
		weights[3846] <= 241;
		weights[3847] <= 3;
		weights[3848] <= 177;
		weights[3849] <= 41;
		weights[3850] <= 54;
		weights[3851] <= 178;
		weights[3852] <= 86;
		weights[3853] <= 132;
		weights[3854] <= 172;
		weights[3855] <= 214;
		weights[3856] <= 205;
		weights[3857] <= 236;
		weights[3858] <= 143;
		weights[3859] <= 231;
		weights[3860] <= 48;
		weights[3861] <= 169;
		weights[3862] <= 231;
		weights[3863] <= 213;
		weights[3864] <= 253;
		weights[3865] <= 8;
		weights[3866] <= 101;
		weights[3867] <= 202;
		weights[3868] <= 131;
		weights[3869] <= 174;
		weights[3870] <= 93;
		weights[3871] <= 95;
		weights[3872] <= 112;
		weights[3873] <= 54;
		weights[3874] <= 233;
		weights[3875] <= 128;
		weights[3876] <= 35;
		weights[3877] <= 152;
		weights[3878] <= 177;
		weights[3879] <= 209;
		weights[3880] <= 32;
		weights[3881] <= 182;
		weights[3882] <= 51;
		weights[3883] <= 150;
		weights[3884] <= 38;
		weights[3885] <= 249;
		weights[3886] <= 115;
		weights[3887] <= 43;
		weights[3888] <= 119;
		weights[3889] <= 38;
		weights[3890] <= 248;
		weights[3891] <= 74;
		weights[3892] <= 90;
		weights[3893] <= 49;
		weights[3894] <= 245;
		weights[3895] <= 227;
		weights[3896] <= 243;
		weights[3897] <= 156;
		weights[3898] <= 94;
		weights[3899] <= 25;
		weights[3900] <= 254;
		weights[3901] <= 72;
		weights[3902] <= 153;
		weights[3903] <= 135;
		weights[3904] <= 97;
		weights[3905] <= 182;
		weights[3906] <= 145;
		weights[3907] <= 173;
		weights[3908] <= 104;
		weights[3909] <= 153;
		weights[3910] <= 101;
		weights[3911] <= 31;
		weights[3912] <= 221;
		weights[3913] <= 192;
		weights[3914] <= 47;
		weights[3915] <= 60;
		weights[3916] <= 123;
		weights[3917] <= 4;
		weights[3918] <= 11;
		weights[3919] <= 60;
		weights[3920] <= 149;
		weights[3921] <= 71;
		weights[3922] <= 159;
		weights[3923] <= 213;
		weights[3924] <= 110;
		weights[3925] <= 18;
		weights[3926] <= 209;
		weights[3927] <= 39;
		weights[3928] <= 190;
		weights[3929] <= 146;
		weights[3930] <= 44;
		weights[3931] <= 88;
		weights[3932] <= 21;
		weights[3933] <= 52;
		weights[3934] <= 93;
		weights[3935] <= 101;
		weights[3936] <= 255;
		weights[3937] <= 100;
		weights[3938] <= 45;
		weights[3939] <= 56;
		weights[3940] <= 107;
		weights[3941] <= 16;
		weights[3942] <= 52;
		weights[3943] <= 77;
		weights[3944] <= 141;
		weights[3945] <= 125;
		weights[3946] <= 125;
		weights[3947] <= 221;
		weights[3948] <= 229;
		weights[3949] <= 4;
		weights[3950] <= 239;
		weights[3951] <= 133;
		weights[3952] <= 245;
		weights[3953] <= 52;
		weights[3954] <= 10;
		weights[3955] <= 30;
		weights[3956] <= 132;
		weights[3957] <= 144;
		weights[3958] <= 21;
		weights[3959] <= 50;
		weights[3960] <= 215;
		weights[3961] <= 160;
		weights[3962] <= 92;
		weights[3963] <= 55;
		weights[3964] <= 124;
		weights[3965] <= 62;
		weights[3966] <= 143;
		weights[3967] <= 142;
		weights[3968] <= 208;
		weights[3969] <= 37;
		weights[3970] <= 38;
		weights[3971] <= 253;
		weights[3972] <= 170;
		weights[3973] <= 240;
		weights[3974] <= 43;
		weights[3975] <= 199;
		weights[3976] <= 79;
		weights[3977] <= 74;
		weights[3978] <= 237;
		weights[3979] <= 80;
		weights[3980] <= 242;
		weights[3981] <= 14;
		weights[3982] <= 126;
		weights[3983] <= 248;
		weights[3984] <= 78;
		weights[3985] <= 44;
		weights[3986] <= 168;
		weights[3987] <= 36;
		weights[3988] <= 201;
		weights[3989] <= 55;
		weights[3990] <= 147;
		weights[3991] <= 3;
		weights[3992] <= 165;
		weights[3993] <= 70;
		weights[3994] <= 3;
		weights[3995] <= 164;
		weights[3996] <= 106;
		weights[3997] <= 72;
		weights[3998] <= 254;
		weights[3999] <= 122;
		weights[4000] <= 26;
		weights[4001] <= 158;
		weights[4002] <= 73;
		weights[4003] <= 15;
		weights[4004] <= 163;
		weights[4005] <= 177;
		weights[4006] <= 67;
		weights[4007] <= 147;
		weights[4008] <= 190;
		weights[4009] <= 246;
		weights[4010] <= 69;
		weights[4011] <= 159;
		weights[4012] <= 221;
		weights[4013] <= 130;
		weights[4014] <= 177;
		weights[4015] <= 114;
		weights[4016] <= 129;
		weights[4017] <= 86;
		weights[4018] <= 199;
		weights[4019] <= 23;
		weights[4020] <= 174;
		weights[4021] <= 176;
		weights[4022] <= 58;
		weights[4023] <= 72;
		weights[4024] <= 50;
		weights[4025] <= 76;
		weights[4026] <= 234;
		weights[4027] <= 195;
		weights[4028] <= 197;
		weights[4029] <= 116;
		weights[4030] <= 204;
		weights[4031] <= 102;
		weights[4032] <= 220;
		weights[4033] <= 220;
		weights[4034] <= 113;
		weights[4035] <= 187;
		weights[4036] <= 16;
		weights[4037] <= 164;
		weights[4038] <= 127;
		weights[4039] <= 238;
		weights[4040] <= 49;
		weights[4041] <= 116;
		weights[4042] <= 194;
		weights[4043] <= 32;
		weights[4044] <= 47;
		weights[4045] <= 65;
		weights[4046] <= 101;
		weights[4047] <= 190;
		weights[4048] <= 154;
		weights[4049] <= 192;
		weights[4050] <= 193;
	end


	always @(negedge(clk)) begin
		if(enable) begin
			case(address)
				12'd0		: data1 <= weights[0];
				12'd1		: data1 <= weights[1];
				12'd2		: data1 <= weights[2];
				12'd3		: data1 <= weights[3];
				12'd4		: data1 <= weights[4];
				12'd5		: data1 <= weights[5];
				12'd6		: data1 <= weights[6];
				12'd7		: data1 <= weights[7];
				12'd8		: data1 <= weights[8];
				12'd9		: data1 <= weights[9];
				12'd10		: data1 <= weights[10];
				12'd11		: data1 <= weights[11];
				12'd12		: data1 <= weights[12];
				12'd13		: data1 <= weights[13];
				12'd14		: data1 <= weights[14];
				12'd15		: data1 <= weights[15];
				12'd16		: data1 <= weights[16];
				12'd17		: data1 <= weights[17];
				12'd18		: data1 <= weights[18];
				12'd19		: data1 <= weights[19];
				12'd20		: data1 <= weights[20];
				12'd21		: data1 <= weights[21];
				12'd22		: data1 <= weights[22];
				12'd23		: data1 <= weights[23];
				12'd24		: data1 <= weights[24];
				12'd25		: data1 <= weights[25];
				12'd26		: data1 <= weights[26];
				12'd27		: data1 <= weights[27];
				12'd28		: data1 <= weights[28];
				12'd29		: data1 <= weights[29];
				12'd30		: data1 <= weights[30];
				12'd31		: data1 <= weights[31];
				12'd32		: data1 <= weights[32];
				12'd33		: data1 <= weights[33];
				12'd34		: data1 <= weights[34];
				12'd35		: data1 <= weights[35];
				12'd36		: data1 <= weights[36];
				12'd37		: data1 <= weights[37];
				12'd38		: data1 <= weights[38];
				12'd39		: data1 <= weights[39];
				12'd40		: data1 <= weights[40];
				12'd41		: data1 <= weights[41];
				12'd42		: data1 <= weights[42];
				12'd43		: data1 <= weights[43];
				12'd44		: data1 <= weights[44];
				12'd45		: data1 <= weights[45];
				12'd46		: data1 <= weights[46];
				12'd47		: data1 <= weights[47];
				12'd48		: data1 <= weights[48];
				12'd49		: data1 <= weights[49];
				12'd50		: data1 <= weights[50];
				12'd51		: data1 <= weights[51];
				12'd52		: data1 <= weights[52];
				12'd53		: data1 <= weights[53];
				12'd54		: data1 <= weights[54];
				12'd55		: data1 <= weights[55];
				12'd56		: data1 <= weights[56];
				12'd57		: data1 <= weights[57];
				12'd58		: data1 <= weights[58];
				12'd59		: data1 <= weights[59];
				12'd60		: data1 <= weights[60];
				12'd61		: data1 <= weights[61];
				12'd62		: data1 <= weights[62];
				12'd63		: data1 <= weights[63];
				12'd64		: data1 <= weights[64];
				12'd65		: data1 <= weights[65];
				12'd66		: data1 <= weights[66];
				12'd67		: data1 <= weights[67];
				12'd68		: data1 <= weights[68];
				12'd69		: data1 <= weights[69];
				12'd70		: data1 <= weights[70];
				12'd71		: data1 <= weights[71];
				12'd72		: data1 <= weights[72];
				12'd73		: data1 <= weights[73];
				12'd74		: data1 <= weights[74];
				12'd75		: data1 <= weights[75];
				12'd76		: data1 <= weights[76];
				12'd77		: data1 <= weights[77];
				12'd78		: data1 <= weights[78];
				12'd79		: data1 <= weights[79];
				12'd80		: data1 <= weights[80];
				12'd81		: data1 <= weights[81];
				12'd82		: data1 <= weights[82];
				12'd83		: data1 <= weights[83];
				12'd84		: data1 <= weights[84];
				12'd85		: data1 <= weights[85];
				12'd86		: data1 <= weights[86];
				12'd87		: data1 <= weights[87];
				12'd88		: data1 <= weights[88];
				12'd89		: data1 <= weights[89];
				12'd90		: data1 <= weights[90];
				12'd91		: data1 <= weights[91];
				12'd92		: data1 <= weights[92];
				12'd93		: data1 <= weights[93];
				12'd94		: data1 <= weights[94];
				12'd95		: data1 <= weights[95];
				12'd96		: data1 <= weights[96];
				12'd97		: data1 <= weights[97];
				12'd98		: data1 <= weights[98];
				12'd99		: data1 <= weights[99];
				12'd100		: data1 <= weights[100];
				12'd101		: data1 <= weights[101];
				12'd102		: data1 <= weights[102];
				12'd103		: data1 <= weights[103];
				12'd104		: data1 <= weights[104];
				12'd105		: data1 <= weights[105];
				12'd106		: data1 <= weights[106];
				12'd107		: data1 <= weights[107];
				12'd108		: data1 <= weights[108];
				12'd109		: data1 <= weights[109];
				12'd110		: data1 <= weights[110];
				12'd111		: data1 <= weights[111];
				12'd112		: data1 <= weights[112];
				12'd113		: data1 <= weights[113];
				12'd114		: data1 <= weights[114];
				12'd115		: data1 <= weights[115];
				12'd116		: data1 <= weights[116];
				12'd117		: data1 <= weights[117];
				12'd118		: data1 <= weights[118];
				12'd119		: data1 <= weights[119];
				12'd120		: data1 <= weights[120];
				12'd121		: data1 <= weights[121];
				12'd122		: data1 <= weights[122];
				12'd123		: data1 <= weights[123];
				12'd124		: data1 <= weights[124];
				12'd125		: data1 <= weights[125];
				12'd126		: data1 <= weights[126];
				12'd127		: data1 <= weights[127];
				12'd128		: data1 <= weights[128];
				12'd129		: data1 <= weights[129];
				12'd130		: data1 <= weights[130];
				12'd131		: data1 <= weights[131];
				12'd132		: data1 <= weights[132];
				12'd133		: data1 <= weights[133];
				12'd134		: data1 <= weights[134];
				12'd135		: data1 <= weights[135];
				12'd136		: data1 <= weights[136];
				12'd137		: data1 <= weights[137];
				12'd138		: data1 <= weights[138];
				12'd139		: data1 <= weights[139];
				12'd140		: data1 <= weights[140];
				12'd141		: data1 <= weights[141];
				12'd142		: data1 <= weights[142];
				12'd143		: data1 <= weights[143];
				12'd144		: data1 <= weights[144];
				12'd145		: data1 <= weights[145];
				12'd146		: data1 <= weights[146];
				12'd147		: data1 <= weights[147];
				12'd148		: data1 <= weights[148];
				12'd149		: data1 <= weights[149];
				12'd150		: data1 <= weights[150];
				12'd151		: data1 <= weights[151];
				12'd152		: data1 <= weights[152];
				12'd153		: data1 <= weights[153];
				12'd154		: data1 <= weights[154];
				12'd155		: data1 <= weights[155];
				12'd156		: data1 <= weights[156];
				12'd157		: data1 <= weights[157];
				12'd158		: data1 <= weights[158];
				12'd159		: data1 <= weights[159];
				12'd160		: data1 <= weights[160];
				12'd161		: data1 <= weights[161];
				12'd162		: data1 <= weights[162];
				12'd163		: data1 <= weights[163];
				12'd164		: data1 <= weights[164];
				12'd165		: data1 <= weights[165];
				12'd166		: data1 <= weights[166];
				12'd167		: data1 <= weights[167];
				12'd168		: data1 <= weights[168];
				12'd169		: data1 <= weights[169];
				12'd170		: data1 <= weights[170];
				12'd171		: data1 <= weights[171];
				12'd172		: data1 <= weights[172];
				12'd173		: data1 <= weights[173];
				12'd174		: data1 <= weights[174];
				12'd175		: data1 <= weights[175];
				12'd176		: data1 <= weights[176];
				12'd177		: data1 <= weights[177];
				12'd178		: data1 <= weights[178];
				12'd179		: data1 <= weights[179];
				12'd180		: data1 <= weights[180];
				12'd181		: data1 <= weights[181];
				12'd182		: data1 <= weights[182];
				12'd183		: data1 <= weights[183];
				12'd184		: data1 <= weights[184];
				12'd185		: data1 <= weights[185];
				12'd186		: data1 <= weights[186];
				12'd187		: data1 <= weights[187];
				12'd188		: data1 <= weights[188];
				12'd189		: data1 <= weights[189];
				12'd190		: data1 <= weights[190];
				12'd191		: data1 <= weights[191];
				12'd192		: data1 <= weights[192];
				12'd193		: data1 <= weights[193];
				12'd194		: data1 <= weights[194];
				12'd195		: data1 <= weights[195];
				12'd196		: data1 <= weights[196];
				12'd197		: data1 <= weights[197];
				12'd198		: data1 <= weights[198];
				12'd199		: data1 <= weights[199];
				12'd200		: data1 <= weights[200];
				12'd201		: data1 <= weights[201];
				12'd202		: data1 <= weights[202];
				12'd203		: data1 <= weights[203];
				12'd204		: data1 <= weights[204];
				12'd205		: data1 <= weights[205];
				12'd206		: data1 <= weights[206];
				12'd207		: data1 <= weights[207];
				12'd208		: data1 <= weights[208];
				12'd209		: data1 <= weights[209];
				12'd210		: data1 <= weights[210];
				12'd211		: data1 <= weights[211];
				12'd212		: data1 <= weights[212];
				12'd213		: data1 <= weights[213];
				12'd214		: data1 <= weights[214];
				12'd215		: data1 <= weights[215];
				12'd216		: data1 <= weights[216];
				12'd217		: data1 <= weights[217];
				12'd218		: data1 <= weights[218];
				12'd219		: data1 <= weights[219];
				12'd220		: data1 <= weights[220];
				12'd221		: data1 <= weights[221];
				12'd222		: data1 <= weights[222];
				12'd223		: data1 <= weights[223];
				12'd224		: data1 <= weights[224];
				12'd225		: data1 <= weights[225];
				12'd226		: data1 <= weights[226];
				12'd227		: data1 <= weights[227];
				12'd228		: data1 <= weights[228];
				12'd229		: data1 <= weights[229];
				12'd230		: data1 <= weights[230];
				12'd231		: data1 <= weights[231];
				12'd232		: data1 <= weights[232];
				12'd233		: data1 <= weights[233];
				12'd234		: data1 <= weights[234];
				12'd235		: data1 <= weights[235];
				12'd236		: data1 <= weights[236];
				12'd237		: data1 <= weights[237];
				12'd238		: data1 <= weights[238];
				12'd239		: data1 <= weights[239];
				12'd240		: data1 <= weights[240];
				12'd241		: data1 <= weights[241];
				12'd242		: data1 <= weights[242];
				12'd243		: data1 <= weights[243];
				12'd244		: data1 <= weights[244];
				12'd245		: data1 <= weights[245];
				12'd246		: data1 <= weights[246];
				12'd247		: data1 <= weights[247];
				12'd248		: data1 <= weights[248];
				12'd249		: data1 <= weights[249];
				12'd250		: data1 <= weights[250];
				12'd251		: data1 <= weights[251];
				12'd252		: data1 <= weights[252];
				12'd253		: data1 <= weights[253];
				12'd254		: data1 <= weights[254];
				12'd255		: data1 <= weights[255];
				12'd256		: data1 <= weights[256];
				12'd257		: data1 <= weights[257];
				12'd258		: data1 <= weights[258];
				12'd259		: data1 <= weights[259];
				12'd260		: data1 <= weights[260];
				12'd261		: data1 <= weights[261];
				12'd262		: data1 <= weights[262];
				12'd263		: data1 <= weights[263];
				12'd264		: data1 <= weights[264];
				12'd265		: data1 <= weights[265];
				12'd266		: data1 <= weights[266];
				12'd267		: data1 <= weights[267];
				12'd268		: data1 <= weights[268];
				12'd269		: data1 <= weights[269];
				12'd270		: data1 <= weights[270];
				12'd271		: data1 <= weights[271];
				12'd272		: data1 <= weights[272];
				12'd273		: data1 <= weights[273];
				12'd274		: data1 <= weights[274];
				12'd275		: data1 <= weights[275];
				12'd276		: data1 <= weights[276];
				12'd277		: data1 <= weights[277];
				12'd278		: data1 <= weights[278];
				12'd279		: data1 <= weights[279];
				12'd280		: data1 <= weights[280];
				12'd281		: data1 <= weights[281];
				12'd282		: data1 <= weights[282];
				12'd283		: data1 <= weights[283];
				12'd284		: data1 <= weights[284];
				12'd285		: data1 <= weights[285];
				12'd286		: data1 <= weights[286];
				12'd287		: data1 <= weights[287];
				12'd288		: data1 <= weights[288];
				12'd289		: data1 <= weights[289];
				12'd290		: data1 <= weights[290];
				12'd291		: data1 <= weights[291];
				12'd292		: data1 <= weights[292];
				12'd293		: data1 <= weights[293];
				12'd294		: data1 <= weights[294];
				12'd295		: data1 <= weights[295];
				12'd296		: data1 <= weights[296];
				12'd297		: data1 <= weights[297];
				12'd298		: data1 <= weights[298];
				12'd299		: data1 <= weights[299];
				12'd300		: data1 <= weights[300];
				12'd301		: data1 <= weights[301];
				12'd302		: data1 <= weights[302];
				12'd303		: data1 <= weights[303];
				12'd304		: data1 <= weights[304];
				12'd305		: data1 <= weights[305];
				12'd306		: data1 <= weights[306];
				12'd307		: data1 <= weights[307];
				12'd308		: data1 <= weights[308];
				12'd309		: data1 <= weights[309];
				12'd310		: data1 <= weights[310];
				12'd311		: data1 <= weights[311];
				12'd312		: data1 <= weights[312];
				12'd313		: data1 <= weights[313];
				12'd314		: data1 <= weights[314];
				12'd315		: data1 <= weights[315];
				12'd316		: data1 <= weights[316];
				12'd317		: data1 <= weights[317];
				12'd318		: data1 <= weights[318];
				12'd319		: data1 <= weights[319];
				12'd320		: data1 <= weights[320];
				12'd321		: data1 <= weights[321];
				12'd322		: data1 <= weights[322];
				12'd323		: data1 <= weights[323];
				12'd324		: data1 <= weights[324];
				12'd325		: data1 <= weights[325];
				12'd326		: data1 <= weights[326];
				12'd327		: data1 <= weights[327];
				12'd328		: data1 <= weights[328];
				12'd329		: data1 <= weights[329];
				12'd330		: data1 <= weights[330];
				12'd331		: data1 <= weights[331];
				12'd332		: data1 <= weights[332];
				12'd333		: data1 <= weights[333];
				12'd334		: data1 <= weights[334];
				12'd335		: data1 <= weights[335];
				12'd336		: data1 <= weights[336];
				12'd337		: data1 <= weights[337];
				12'd338		: data1 <= weights[338];
				12'd339		: data1 <= weights[339];
				12'd340		: data1 <= weights[340];
				12'd341		: data1 <= weights[341];
				12'd342		: data1 <= weights[342];
				12'd343		: data1 <= weights[343];
				12'd344		: data1 <= weights[344];
				12'd345		: data1 <= weights[345];
				12'd346		: data1 <= weights[346];
				12'd347		: data1 <= weights[347];
				12'd348		: data1 <= weights[348];
				12'd349		: data1 <= weights[349];
				12'd350		: data1 <= weights[350];
				12'd351		: data1 <= weights[351];
				12'd352		: data1 <= weights[352];
				12'd353		: data1 <= weights[353];
				12'd354		: data1 <= weights[354];
				12'd355		: data1 <= weights[355];
				12'd356		: data1 <= weights[356];
				12'd357		: data1 <= weights[357];
				12'd358		: data1 <= weights[358];
				12'd359		: data1 <= weights[359];
				12'd360		: data1 <= weights[360];
				12'd361		: data1 <= weights[361];
				12'd362		: data1 <= weights[362];
				12'd363		: data1 <= weights[363];
				12'd364		: data1 <= weights[364];
				12'd365		: data1 <= weights[365];
				12'd366		: data1 <= weights[366];
				12'd367		: data1 <= weights[367];
				12'd368		: data1 <= weights[368];
				12'd369		: data1 <= weights[369];
				12'd370		: data1 <= weights[370];
				12'd371		: data1 <= weights[371];
				12'd372		: data1 <= weights[372];
				12'd373		: data1 <= weights[373];
				12'd374		: data1 <= weights[374];
				12'd375		: data1 <= weights[375];
				12'd376		: data1 <= weights[376];
				12'd377		: data1 <= weights[377];
				12'd378		: data1 <= weights[378];
				12'd379		: data1 <= weights[379];
				12'd380		: data1 <= weights[380];
				12'd381		: data1 <= weights[381];
				12'd382		: data1 <= weights[382];
				12'd383		: data1 <= weights[383];
				12'd384		: data1 <= weights[384];
				12'd385		: data1 <= weights[385];
				12'd386		: data1 <= weights[386];
				12'd387		: data1 <= weights[387];
				12'd388		: data1 <= weights[388];
				12'd389		: data1 <= weights[389];
				12'd390		: data1 <= weights[390];
				12'd391		: data1 <= weights[391];
				12'd392		: data1 <= weights[392];
				12'd393		: data1 <= weights[393];
				12'd394		: data1 <= weights[394];
				12'd395		: data1 <= weights[395];
				12'd396		: data1 <= weights[396];
				12'd397		: data1 <= weights[397];
				12'd398		: data1 <= weights[398];
				12'd399		: data1 <= weights[399];
				12'd400		: data1 <= weights[400];
				12'd401		: data1 <= weights[401];
				12'd402		: data1 <= weights[402];
				12'd403		: data1 <= weights[403];
				12'd404		: data1 <= weights[404];
				12'd405		: data1 <= weights[405];
				12'd406		: data1 <= weights[406];
				12'd407		: data1 <= weights[407];
				12'd408		: data1 <= weights[408];
				12'd409		: data1 <= weights[409];
				12'd410		: data1 <= weights[410];
				12'd411		: data1 <= weights[411];
				12'd412		: data1 <= weights[412];
				12'd413		: data1 <= weights[413];
				12'd414		: data1 <= weights[414];
				12'd415		: data1 <= weights[415];
				12'd416		: data1 <= weights[416];
				12'd417		: data1 <= weights[417];
				12'd418		: data1 <= weights[418];
				12'd419		: data1 <= weights[419];
				12'd420		: data1 <= weights[420];
				12'd421		: data1 <= weights[421];
				12'd422		: data1 <= weights[422];
				12'd423		: data1 <= weights[423];
				12'd424		: data1 <= weights[424];
				12'd425		: data1 <= weights[425];
				12'd426		: data1 <= weights[426];
				12'd427		: data1 <= weights[427];
				12'd428		: data1 <= weights[428];
				12'd429		: data1 <= weights[429];
				12'd430		: data1 <= weights[430];
				12'd431		: data1 <= weights[431];
				12'd432		: data1 <= weights[432];
				12'd433		: data1 <= weights[433];
				12'd434		: data1 <= weights[434];
				12'd435		: data1 <= weights[435];
				12'd436		: data1 <= weights[436];
				12'd437		: data1 <= weights[437];
				12'd438		: data1 <= weights[438];
				12'd439		: data1 <= weights[439];
				12'd440		: data1 <= weights[440];
				12'd441		: data1 <= weights[441];
				12'd442		: data1 <= weights[442];
				12'd443		: data1 <= weights[443];
				12'd444		: data1 <= weights[444];
				12'd445		: data1 <= weights[445];
				12'd446		: data1 <= weights[446];
				12'd447		: data1 <= weights[447];
				12'd448		: data1 <= weights[448];
				12'd449		: data1 <= weights[449];
				12'd450		: data1 <= weights[450];
				12'd451		: data1 <= weights[451];
				12'd452		: data1 <= weights[452];
				12'd453		: data1 <= weights[453];
				12'd454		: data1 <= weights[454];
				12'd455		: data1 <= weights[455];
				12'd456		: data1 <= weights[456];
				12'd457		: data1 <= weights[457];
				12'd458		: data1 <= weights[458];
				12'd459		: data1 <= weights[459];
				12'd460		: data1 <= weights[460];
				12'd461		: data1 <= weights[461];
				12'd462		: data1 <= weights[462];
				12'd463		: data1 <= weights[463];
				12'd464		: data1 <= weights[464];
				12'd465		: data1 <= weights[465];
				12'd466		: data1 <= weights[466];
				12'd467		: data1 <= weights[467];
				12'd468		: data1 <= weights[468];
				12'd469		: data1 <= weights[469];
				12'd470		: data1 <= weights[470];
				12'd471		: data1 <= weights[471];
				12'd472		: data1 <= weights[472];
				12'd473		: data1 <= weights[473];
				12'd474		: data1 <= weights[474];
				12'd475		: data1 <= weights[475];
				12'd476		: data1 <= weights[476];
				12'd477		: data1 <= weights[477];
				12'd478		: data1 <= weights[478];
				12'd479		: data1 <= weights[479];
				12'd480		: data1 <= weights[480];
				12'd481		: data1 <= weights[481];
				12'd482		: data1 <= weights[482];
				12'd483		: data1 <= weights[483];
				12'd484		: data1 <= weights[484];
				12'd485		: data1 <= weights[485];
				12'd486		: data1 <= weights[486];
				12'd487		: data1 <= weights[487];
				12'd488		: data1 <= weights[488];
				12'd489		: data1 <= weights[489];
				12'd490		: data1 <= weights[490];
				12'd491		: data1 <= weights[491];
				12'd492		: data1 <= weights[492];
				12'd493		: data1 <= weights[493];
				12'd494		: data1 <= weights[494];
				12'd495		: data1 <= weights[495];
				12'd496		: data1 <= weights[496];
				12'd497		: data1 <= weights[497];
				12'd498		: data1 <= weights[498];
				12'd499		: data1 <= weights[499];
				12'd500		: data1 <= weights[500];
				12'd501		: data1 <= weights[501];
				12'd502		: data1 <= weights[502];
				12'd503		: data1 <= weights[503];
				12'd504		: data1 <= weights[504];
				12'd505		: data1 <= weights[505];
				12'd506		: data1 <= weights[506];
				12'd507		: data1 <= weights[507];
				12'd508		: data1 <= weights[508];
				12'd509		: data1 <= weights[509];
				12'd510		: data1 <= weights[510];
				12'd511		: data1 <= weights[511];
				12'd512		: data1 <= weights[512];
				12'd513		: data1 <= weights[513];
				12'd514		: data1 <= weights[514];
				12'd515		: data1 <= weights[515];
				12'd516		: data1 <= weights[516];
				12'd517		: data1 <= weights[517];
				12'd518		: data1 <= weights[518];
				12'd519		: data1 <= weights[519];
				12'd520		: data1 <= weights[520];
				12'd521		: data1 <= weights[521];
				12'd522		: data1 <= weights[522];
				12'd523		: data1 <= weights[523];
				12'd524		: data1 <= weights[524];
				12'd525		: data1 <= weights[525];
				12'd526		: data1 <= weights[526];
				12'd527		: data1 <= weights[527];
				12'd528		: data1 <= weights[528];
				12'd529		: data1 <= weights[529];
				12'd530		: data1 <= weights[530];
				12'd531		: data1 <= weights[531];
				12'd532		: data1 <= weights[532];
				12'd533		: data1 <= weights[533];
				12'd534		: data1 <= weights[534];
				12'd535		: data1 <= weights[535];
				12'd536		: data1 <= weights[536];
				12'd537		: data1 <= weights[537];
				12'd538		: data1 <= weights[538];
				12'd539		: data1 <= weights[539];
				12'd540		: data1 <= weights[540];
				12'd541		: data1 <= weights[541];
				12'd542		: data1 <= weights[542];
				12'd543		: data1 <= weights[543];
				12'd544		: data1 <= weights[544];
				12'd545		: data1 <= weights[545];
				12'd546		: data1 <= weights[546];
				12'd547		: data1 <= weights[547];
				12'd548		: data1 <= weights[548];
				12'd549		: data1 <= weights[549];
				12'd550		: data1 <= weights[550];
				12'd551		: data1 <= weights[551];
				12'd552		: data1 <= weights[552];
				12'd553		: data1 <= weights[553];
				12'd554		: data1 <= weights[554];
				12'd555		: data1 <= weights[555];
				12'd556		: data1 <= weights[556];
				12'd557		: data1 <= weights[557];
				12'd558		: data1 <= weights[558];
				12'd559		: data1 <= weights[559];
				12'd560		: data1 <= weights[560];
				12'd561		: data1 <= weights[561];
				12'd562		: data1 <= weights[562];
				12'd563		: data1 <= weights[563];
				12'd564		: data1 <= weights[564];
				12'd565		: data1 <= weights[565];
				12'd566		: data1 <= weights[566];
				12'd567		: data1 <= weights[567];
				12'd568		: data1 <= weights[568];
				12'd569		: data1 <= weights[569];
				12'd570		: data1 <= weights[570];
				12'd571		: data1 <= weights[571];
				12'd572		: data1 <= weights[572];
				12'd573		: data1 <= weights[573];
				12'd574		: data1 <= weights[574];
				12'd575		: data1 <= weights[575];
				12'd576		: data1 <= weights[576];
				12'd577		: data1 <= weights[577];
				12'd578		: data1 <= weights[578];
				12'd579		: data1 <= weights[579];
				12'd580		: data1 <= weights[580];
				12'd581		: data1 <= weights[581];
				12'd582		: data1 <= weights[582];
				12'd583		: data1 <= weights[583];
				12'd584		: data1 <= weights[584];
				12'd585		: data1 <= weights[585];
				12'd586		: data1 <= weights[586];
				12'd587		: data1 <= weights[587];
				12'd588		: data1 <= weights[588];
				12'd589		: data1 <= weights[589];
				12'd590		: data1 <= weights[590];
				12'd591		: data1 <= weights[591];
				12'd592		: data1 <= weights[592];
				12'd593		: data1 <= weights[593];
				12'd594		: data1 <= weights[594];
				12'd595		: data1 <= weights[595];
				12'd596		: data1 <= weights[596];
				12'd597		: data1 <= weights[597];
				12'd598		: data1 <= weights[598];
				12'd599		: data1 <= weights[599];
				12'd600		: data1 <= weights[600];
				12'd601		: data1 <= weights[601];
				12'd602		: data1 <= weights[602];
				12'd603		: data1 <= weights[603];
				12'd604		: data1 <= weights[604];
				12'd605		: data1 <= weights[605];
				12'd606		: data1 <= weights[606];
				12'd607		: data1 <= weights[607];
				12'd608		: data1 <= weights[608];
				12'd609		: data1 <= weights[609];
				12'd610		: data1 <= weights[610];
				12'd611		: data1 <= weights[611];
				12'd612		: data1 <= weights[612];
				12'd613		: data1 <= weights[613];
				12'd614		: data1 <= weights[614];
				12'd615		: data1 <= weights[615];
				12'd616		: data1 <= weights[616];
				12'd617		: data1 <= weights[617];
				12'd618		: data1 <= weights[618];
				12'd619		: data1 <= weights[619];
				12'd620		: data1 <= weights[620];
				12'd621		: data1 <= weights[621];
				12'd622		: data1 <= weights[622];
				12'd623		: data1 <= weights[623];
				12'd624		: data1 <= weights[624];
				12'd625		: data1 <= weights[625];
				12'd626		: data1 <= weights[626];
				12'd627		: data1 <= weights[627];
				12'd628		: data1 <= weights[628];
				12'd629		: data1 <= weights[629];
				12'd630		: data1 <= weights[630];
				12'd631		: data1 <= weights[631];
				12'd632		: data1 <= weights[632];
				12'd633		: data1 <= weights[633];
				12'd634		: data1 <= weights[634];
				12'd635		: data1 <= weights[635];
				12'd636		: data1 <= weights[636];
				12'd637		: data1 <= weights[637];
				12'd638		: data1 <= weights[638];
				12'd639		: data1 <= weights[639];
				12'd640		: data1 <= weights[640];
				12'd641		: data1 <= weights[641];
				12'd642		: data1 <= weights[642];
				12'd643		: data1 <= weights[643];
				12'd644		: data1 <= weights[644];
				12'd645		: data1 <= weights[645];
				12'd646		: data1 <= weights[646];
				12'd647		: data1 <= weights[647];
				12'd648		: data1 <= weights[648];
				12'd649		: data1 <= weights[649];
				12'd650		: data1 <= weights[650];
				12'd651		: data1 <= weights[651];
				12'd652		: data1 <= weights[652];
				12'd653		: data1 <= weights[653];
				12'd654		: data1 <= weights[654];
				12'd655		: data1 <= weights[655];
				12'd656		: data1 <= weights[656];
				12'd657		: data1 <= weights[657];
				12'd658		: data1 <= weights[658];
				12'd659		: data1 <= weights[659];
				12'd660		: data1 <= weights[660];
				12'd661		: data1 <= weights[661];
				12'd662		: data1 <= weights[662];
				12'd663		: data1 <= weights[663];
				12'd664		: data1 <= weights[664];
				12'd665		: data1 <= weights[665];
				12'd666		: data1 <= weights[666];
				12'd667		: data1 <= weights[667];
				12'd668		: data1 <= weights[668];
				12'd669		: data1 <= weights[669];
				12'd670		: data1 <= weights[670];
				12'd671		: data1 <= weights[671];
				12'd672		: data1 <= weights[672];
				12'd673		: data1 <= weights[673];
				12'd674		: data1 <= weights[674];
				12'd675		: data1 <= weights[675];
				12'd676		: data1 <= weights[676];
				12'd677		: data1 <= weights[677];
				12'd678		: data1 <= weights[678];
				12'd679		: data1 <= weights[679];
				12'd680		: data1 <= weights[680];
				12'd681		: data1 <= weights[681];
				12'd682		: data1 <= weights[682];
				12'd683		: data1 <= weights[683];
				12'd684		: data1 <= weights[684];
				12'd685		: data1 <= weights[685];
				12'd686		: data1 <= weights[686];
				12'd687		: data1 <= weights[687];
				12'd688		: data1 <= weights[688];
				12'd689		: data1 <= weights[689];
				12'd690		: data1 <= weights[690];
				12'd691		: data1 <= weights[691];
				12'd692		: data1 <= weights[692];
				12'd693		: data1 <= weights[693];
				12'd694		: data1 <= weights[694];
				12'd695		: data1 <= weights[695];
				12'd696		: data1 <= weights[696];
				12'd697		: data1 <= weights[697];
				12'd698		: data1 <= weights[698];
				12'd699		: data1 <= weights[699];
				12'd700		: data1 <= weights[700];
				12'd701		: data1 <= weights[701];
				12'd702		: data1 <= weights[702];
				12'd703		: data1 <= weights[703];
				12'd704		: data1 <= weights[704];
				12'd705		: data1 <= weights[705];
				12'd706		: data1 <= weights[706];
				12'd707		: data1 <= weights[707];
				12'd708		: data1 <= weights[708];
				12'd709		: data1 <= weights[709];
				12'd710		: data1 <= weights[710];
				12'd711		: data1 <= weights[711];
				12'd712		: data1 <= weights[712];
				12'd713		: data1 <= weights[713];
				12'd714		: data1 <= weights[714];
				12'd715		: data1 <= weights[715];
				12'd716		: data1 <= weights[716];
				12'd717		: data1 <= weights[717];
				12'd718		: data1 <= weights[718];
				12'd719		: data1 <= weights[719];
				12'd720		: data1 <= weights[720];
				12'd721		: data1 <= weights[721];
				12'd722		: data1 <= weights[722];
				12'd723		: data1 <= weights[723];
				12'd724		: data1 <= weights[724];
				12'd725		: data1 <= weights[725];
				12'd726		: data1 <= weights[726];
				12'd727		: data1 <= weights[727];
				12'd728		: data1 <= weights[728];
				12'd729		: data1 <= weights[729];
				12'd730		: data1 <= weights[730];
				12'd731		: data1 <= weights[731];
				12'd732		: data1 <= weights[732];
				12'd733		: data1 <= weights[733];
				12'd734		: data1 <= weights[734];
				12'd735		: data1 <= weights[735];
				12'd736		: data1 <= weights[736];
				12'd737		: data1 <= weights[737];
				12'd738		: data1 <= weights[738];
				12'd739		: data1 <= weights[739];
				12'd740		: data1 <= weights[740];
				12'd741		: data1 <= weights[741];
				12'd742		: data1 <= weights[742];
				12'd743		: data1 <= weights[743];
				12'd744		: data1 <= weights[744];
				12'd745		: data1 <= weights[745];
				12'd746		: data1 <= weights[746];
				12'd747		: data1 <= weights[747];
				12'd748		: data1 <= weights[748];
				12'd749		: data1 <= weights[749];
				12'd750		: data1 <= weights[750];
				12'd751		: data1 <= weights[751];
				12'd752		: data1 <= weights[752];
				12'd753		: data1 <= weights[753];
				12'd754		: data1 <= weights[754];
				12'd755		: data1 <= weights[755];
				12'd756		: data1 <= weights[756];
				12'd757		: data1 <= weights[757];
				12'd758		: data1 <= weights[758];
				12'd759		: data1 <= weights[759];
				12'd760		: data1 <= weights[760];
				12'd761		: data1 <= weights[761];
				12'd762		: data1 <= weights[762];
				12'd763		: data1 <= weights[763];
				12'd764		: data1 <= weights[764];
				12'd765		: data1 <= weights[765];
				12'd766		: data1 <= weights[766];
				12'd767		: data1 <= weights[767];
				12'd768		: data1 <= weights[768];
				12'd769		: data1 <= weights[769];
				12'd770		: data1 <= weights[770];
				12'd771		: data1 <= weights[771];
				12'd772		: data1 <= weights[772];
				12'd773		: data1 <= weights[773];
				12'd774		: data1 <= weights[774];
				12'd775		: data1 <= weights[775];
				12'd776		: data1 <= weights[776];
				12'd777		: data1 <= weights[777];
				12'd778		: data1 <= weights[778];
				12'd779		: data1 <= weights[779];
				12'd780		: data1 <= weights[780];
				12'd781		: data1 <= weights[781];
				12'd782		: data1 <= weights[782];
				12'd783		: data1 <= weights[783];
				12'd784		: data1 <= weights[784];
				12'd785		: data1 <= weights[785];
				12'd786		: data1 <= weights[786];
				12'd787		: data1 <= weights[787];
				12'd788		: data1 <= weights[788];
				12'd789		: data1 <= weights[789];
				12'd790		: data1 <= weights[790];
				12'd791		: data1 <= weights[791];
				12'd792		: data1 <= weights[792];
				12'd793		: data1 <= weights[793];
				12'd794		: data1 <= weights[794];
				12'd795		: data1 <= weights[795];
				12'd796		: data1 <= weights[796];
				12'd797		: data1 <= weights[797];
				12'd798		: data1 <= weights[798];
				12'd799		: data1 <= weights[799];
				12'd800		: data1 <= weights[800];
				12'd801		: data1 <= weights[801];
				12'd802		: data1 <= weights[802];
				12'd803		: data1 <= weights[803];
				12'd804		: data1 <= weights[804];
				12'd805		: data1 <= weights[805];
				12'd806		: data1 <= weights[806];
				12'd807		: data1 <= weights[807];
				12'd808		: data1 <= weights[808];
				12'd809		: data1 <= weights[809];
				12'd810		: data1 <= weights[810];
				12'd811		: data1 <= weights[811];
				12'd812		: data1 <= weights[812];
				12'd813		: data1 <= weights[813];
				12'd814		: data1 <= weights[814];
				12'd815		: data1 <= weights[815];
				12'd816		: data1 <= weights[816];
				12'd817		: data1 <= weights[817];
				12'd818		: data1 <= weights[818];
				12'd819		: data1 <= weights[819];
				12'd820		: data1 <= weights[820];
				12'd821		: data1 <= weights[821];
				12'd822		: data1 <= weights[822];
				12'd823		: data1 <= weights[823];
				12'd824		: data1 <= weights[824];
				12'd825		: data1 <= weights[825];
				12'd826		: data1 <= weights[826];
				12'd827		: data1 <= weights[827];
				12'd828		: data1 <= weights[828];
				12'd829		: data1 <= weights[829];
				12'd830		: data1 <= weights[830];
				12'd831		: data1 <= weights[831];
				12'd832		: data1 <= weights[832];
				12'd833		: data1 <= weights[833];
				12'd834		: data1 <= weights[834];
				12'd835		: data1 <= weights[835];
				12'd836		: data1 <= weights[836];
				12'd837		: data1 <= weights[837];
				12'd838		: data1 <= weights[838];
				12'd839		: data1 <= weights[839];
				12'd840		: data1 <= weights[840];
				12'd841		: data1 <= weights[841];
				12'd842		: data1 <= weights[842];
				12'd843		: data1 <= weights[843];
				12'd844		: data1 <= weights[844];
				12'd845		: data1 <= weights[845];
				12'd846		: data1 <= weights[846];
				12'd847		: data1 <= weights[847];
				12'd848		: data1 <= weights[848];
				12'd849		: data1 <= weights[849];
				12'd850		: data1 <= weights[850];
				12'd851		: data1 <= weights[851];
				12'd852		: data1 <= weights[852];
				12'd853		: data1 <= weights[853];
				12'd854		: data1 <= weights[854];
				12'd855		: data1 <= weights[855];
				12'd856		: data1 <= weights[856];
				12'd857		: data1 <= weights[857];
				12'd858		: data1 <= weights[858];
				12'd859		: data1 <= weights[859];
				12'd860		: data1 <= weights[860];
				12'd861		: data1 <= weights[861];
				12'd862		: data1 <= weights[862];
				12'd863		: data1 <= weights[863];
				12'd864		: data1 <= weights[864];
				12'd865		: data1 <= weights[865];
				12'd866		: data1 <= weights[866];
				12'd867		: data1 <= weights[867];
				12'd868		: data1 <= weights[868];
				12'd869		: data1 <= weights[869];
				12'd870		: data1 <= weights[870];
				12'd871		: data1 <= weights[871];
				12'd872		: data1 <= weights[872];
				12'd873		: data1 <= weights[873];
				12'd874		: data1 <= weights[874];
				12'd875		: data1 <= weights[875];
				12'd876		: data1 <= weights[876];
				12'd877		: data1 <= weights[877];
				12'd878		: data1 <= weights[878];
				12'd879		: data1 <= weights[879];
				12'd880		: data1 <= weights[880];
				12'd881		: data1 <= weights[881];
				12'd882		: data1 <= weights[882];
				12'd883		: data1 <= weights[883];
				12'd884		: data1 <= weights[884];
				12'd885		: data1 <= weights[885];
				12'd886		: data1 <= weights[886];
				12'd887		: data1 <= weights[887];
				12'd888		: data1 <= weights[888];
				12'd889		: data1 <= weights[889];
				12'd890		: data1 <= weights[890];
				12'd891		: data1 <= weights[891];
				12'd892		: data1 <= weights[892];
				12'd893		: data1 <= weights[893];
				12'd894		: data1 <= weights[894];
				12'd895		: data1 <= weights[895];
				12'd896		: data1 <= weights[896];
				12'd897		: data1 <= weights[897];
				12'd898		: data1 <= weights[898];
				12'd899		: data1 <= weights[899];
				12'd900		: data1 <= weights[900];
				12'd901		: data1 <= weights[901];
				12'd902		: data1 <= weights[902];
				12'd903		: data1 <= weights[903];
				12'd904		: data1 <= weights[904];
				12'd905		: data1 <= weights[905];
				12'd906		: data1 <= weights[906];
				12'd907		: data1 <= weights[907];
				12'd908		: data1 <= weights[908];
				12'd909		: data1 <= weights[909];
				12'd910		: data1 <= weights[910];
				12'd911		: data1 <= weights[911];
				12'd912		: data1 <= weights[912];
				12'd913		: data1 <= weights[913];
				12'd914		: data1 <= weights[914];
				12'd915		: data1 <= weights[915];
				12'd916		: data1 <= weights[916];
				12'd917		: data1 <= weights[917];
				12'd918		: data1 <= weights[918];
				12'd919		: data1 <= weights[919];
				12'd920		: data1 <= weights[920];
				12'd921		: data1 <= weights[921];
				12'd922		: data1 <= weights[922];
				12'd923		: data1 <= weights[923];
				12'd924		: data1 <= weights[924];
				12'd925		: data1 <= weights[925];
				12'd926		: data1 <= weights[926];
				12'd927		: data1 <= weights[927];
				12'd928		: data1 <= weights[928];
				12'd929		: data1 <= weights[929];
				12'd930		: data1 <= weights[930];
				12'd931		: data1 <= weights[931];
				12'd932		: data1 <= weights[932];
				12'd933		: data1 <= weights[933];
				12'd934		: data1 <= weights[934];
				12'd935		: data1 <= weights[935];
				12'd936		: data1 <= weights[936];
				12'd937		: data1 <= weights[937];
				12'd938		: data1 <= weights[938];
				12'd939		: data1 <= weights[939];
				12'd940		: data1 <= weights[940];
				12'd941		: data1 <= weights[941];
				12'd942		: data1 <= weights[942];
				12'd943		: data1 <= weights[943];
				12'd944		: data1 <= weights[944];
				12'd945		: data1 <= weights[945];
				12'd946		: data1 <= weights[946];
				12'd947		: data1 <= weights[947];
				12'd948		: data1 <= weights[948];
				12'd949		: data1 <= weights[949];
				12'd950		: data1 <= weights[950];
				12'd951		: data1 <= weights[951];
				12'd952		: data1 <= weights[952];
				12'd953		: data1 <= weights[953];
				12'd954		: data1 <= weights[954];
				12'd955		: data1 <= weights[955];
				12'd956		: data1 <= weights[956];
				12'd957		: data1 <= weights[957];
				12'd958		: data1 <= weights[958];
				12'd959		: data1 <= weights[959];
				12'd960		: data1 <= weights[960];
				12'd961		: data1 <= weights[961];
				12'd962		: data1 <= weights[962];
				12'd963		: data1 <= weights[963];
				12'd964		: data1 <= weights[964];
				12'd965		: data1 <= weights[965];
				12'd966		: data1 <= weights[966];
				12'd967		: data1 <= weights[967];
				12'd968		: data1 <= weights[968];
				12'd969		: data1 <= weights[969];
				12'd970		: data1 <= weights[970];
				12'd971		: data1 <= weights[971];
				12'd972		: data1 <= weights[972];
				12'd973		: data1 <= weights[973];
				12'd974		: data1 <= weights[974];
				12'd975		: data1 <= weights[975];
				12'd976		: data1 <= weights[976];
				12'd977		: data1 <= weights[977];
				12'd978		: data1 <= weights[978];
				12'd979		: data1 <= weights[979];
				12'd980		: data1 <= weights[980];
				12'd981		: data1 <= weights[981];
				12'd982		: data1 <= weights[982];
				12'd983		: data1 <= weights[983];
				12'd984		: data1 <= weights[984];
				12'd985		: data1 <= weights[985];
				12'd986		: data1 <= weights[986];
				12'd987		: data1 <= weights[987];
				12'd988		: data1 <= weights[988];
				12'd989		: data1 <= weights[989];
				12'd990		: data1 <= weights[990];
				12'd991		: data1 <= weights[991];
				12'd992		: data1 <= weights[992];
				12'd993		: data1 <= weights[993];
				12'd994		: data1 <= weights[994];
				12'd995		: data1 <= weights[995];
				12'd996		: data1 <= weights[996];
				12'd997		: data1 <= weights[997];
				12'd998		: data1 <= weights[998];
				12'd999		: data1 <= weights[999];
				12'd1000	: data1 <= weights[1000];
				12'd1001	: data1 <= weights[1001];
				12'd1002	: data1 <= weights[1002];
				12'd1003	: data1 <= weights[1003];
				12'd1004	: data1 <= weights[1004];
				12'd1005	: data1 <= weights[1005];
				12'd1006	: data1 <= weights[1006];
				12'd1007	: data1 <= weights[1007];
				12'd1008	: data1 <= weights[1008];
				12'd1009	: data1 <= weights[1009];
				12'd1010	: data1 <= weights[1010];
				12'd1011	: data1 <= weights[1011];
				12'd1012	: data1 <= weights[1012];
				12'd1013	: data1 <= weights[1013];
				12'd1014	: data1 <= weights[1014];
				12'd1015	: data1 <= weights[1015];
				12'd1016	: data1 <= weights[1016];
				12'd1017	: data1 <= weights[1017];
				12'd1018	: data1 <= weights[1018];
				12'd1019	: data1 <= weights[1019];
				12'd1020	: data1 <= weights[1020];
				12'd1021	: data1 <= weights[1021];
				12'd1022	: data1 <= weights[1022];
				12'd1023	: data1 <= weights[1023];
				12'd1024	: data1 <= weights[1024];
				12'd1025	: data1 <= weights[1025];
				12'd1026	: data1 <= weights[1026];
				12'd1027	: data1 <= weights[1027];
				12'd1028	: data1 <= weights[1028];
				12'd1029	: data1 <= weights[1029];
				12'd1030	: data1 <= weights[1030];
				12'd1031	: data1 <= weights[1031];
				12'd1032	: data1 <= weights[1032];
				12'd1033	: data1 <= weights[1033];
				12'd1034	: data1 <= weights[1034];
				12'd1035	: data1 <= weights[1035];
				12'd1036	: data1 <= weights[1036];
				12'd1037	: data1 <= weights[1037];
				12'd1038	: data1 <= weights[1038];
				12'd1039	: data1 <= weights[1039];
				12'd1040	: data1 <= weights[1040];
				12'd1041	: data1 <= weights[1041];
				12'd1042	: data1 <= weights[1042];
				12'd1043	: data1 <= weights[1043];
				12'd1044	: data1 <= weights[1044];
				12'd1045	: data1 <= weights[1045];
				12'd1046	: data1 <= weights[1046];
				12'd1047	: data1 <= weights[1047];
				12'd1048	: data1 <= weights[1048];
				12'd1049	: data1 <= weights[1049];
				12'd1050	: data1 <= weights[1050];
				12'd1051	: data1 <= weights[1051];
				12'd1052	: data1 <= weights[1052];
				12'd1053	: data1 <= weights[1053];
				12'd1054	: data1 <= weights[1054];
				12'd1055	: data1 <= weights[1055];
				12'd1056	: data1 <= weights[1056];
				12'd1057	: data1 <= weights[1057];
				12'd1058	: data1 <= weights[1058];
				12'd1059	: data1 <= weights[1059];
				12'd1060	: data1 <= weights[1060];
				12'd1061	: data1 <= weights[1061];
				12'd1062	: data1 <= weights[1062];
				12'd1063	: data1 <= weights[1063];
				12'd1064	: data1 <= weights[1064];
				12'd1065	: data1 <= weights[1065];
				12'd1066	: data1 <= weights[1066];
				12'd1067	: data1 <= weights[1067];
				12'd1068	: data1 <= weights[1068];
				12'd1069	: data1 <= weights[1069];
				12'd1070	: data1 <= weights[1070];
				12'd1071	: data1 <= weights[1071];
				12'd1072	: data1 <= weights[1072];
				12'd1073	: data1 <= weights[1073];
				12'd1074	: data1 <= weights[1074];
				12'd1075	: data1 <= weights[1075];
				12'd1076	: data1 <= weights[1076];
				12'd1077	: data1 <= weights[1077];
				12'd1078	: data1 <= weights[1078];
				12'd1079	: data1 <= weights[1079];
				12'd1080	: data1 <= weights[1080];
				12'd1081	: data1 <= weights[1081];
				12'd1082	: data1 <= weights[1082];
				12'd1083	: data1 <= weights[1083];
				12'd1084	: data1 <= weights[1084];
				12'd1085	: data1 <= weights[1085];
				12'd1086	: data1 <= weights[1086];
				12'd1087	: data1 <= weights[1087];
				12'd1088	: data1 <= weights[1088];
				12'd1089	: data1 <= weights[1089];
				12'd1090	: data1 <= weights[1090];
				12'd1091	: data1 <= weights[1091];
				12'd1092	: data1 <= weights[1092];
				12'd1093	: data1 <= weights[1093];
				12'd1094	: data1 <= weights[1094];
				12'd1095	: data1 <= weights[1095];
				12'd1096	: data1 <= weights[1096];
				12'd1097	: data1 <= weights[1097];
				12'd1098	: data1 <= weights[1098];
				12'd1099	: data1 <= weights[1099];
				12'd1100	: data1 <= weights[1100];
				12'd1101	: data1 <= weights[1101];
				12'd1102	: data1 <= weights[1102];
				12'd1103	: data1 <= weights[1103];
				12'd1104	: data1 <= weights[1104];
				12'd1105	: data1 <= weights[1105];
				12'd1106	: data1 <= weights[1106];
				12'd1107	: data1 <= weights[1107];
				12'd1108	: data1 <= weights[1108];
				12'd1109	: data1 <= weights[1109];
				12'd1110	: data1 <= weights[1110];
				12'd1111	: data1 <= weights[1111];
				12'd1112	: data1 <= weights[1112];
				12'd1113	: data1 <= weights[1113];
				12'd1114	: data1 <= weights[1114];
				12'd1115	: data1 <= weights[1115];
				12'd1116	: data1 <= weights[1116];
				12'd1117	: data1 <= weights[1117];
				12'd1118	: data1 <= weights[1118];
				12'd1119	: data1 <= weights[1119];
				12'd1120	: data1 <= weights[1120];
				12'd1121	: data1 <= weights[1121];
				12'd1122	: data1 <= weights[1122];
				12'd1123	: data1 <= weights[1123];
				12'd1124	: data1 <= weights[1124];
				12'd1125	: data1 <= weights[1125];
				12'd1126	: data1 <= weights[1126];
				12'd1127	: data1 <= weights[1127];
				12'd1128	: data1 <= weights[1128];
				12'd1129	: data1 <= weights[1129];
				12'd1130	: data1 <= weights[1130];
				12'd1131	: data1 <= weights[1131];
				12'd1132	: data1 <= weights[1132];
				12'd1133	: data1 <= weights[1133];
				12'd1134	: data1 <= weights[1134];
				12'd1135	: data1 <= weights[1135];
				12'd1136	: data1 <= weights[1136];
				12'd1137	: data1 <= weights[1137];
				12'd1138	: data1 <= weights[1138];
				12'd1139	: data1 <= weights[1139];
				12'd1140	: data1 <= weights[1140];
				12'd1141	: data1 <= weights[1141];
				12'd1142	: data1 <= weights[1142];
				12'd1143	: data1 <= weights[1143];
				12'd1144	: data1 <= weights[1144];
				12'd1145	: data1 <= weights[1145];
				12'd1146	: data1 <= weights[1146];
				12'd1147	: data1 <= weights[1147];
				12'd1148	: data1 <= weights[1148];
				12'd1149	: data1 <= weights[1149];
				12'd1150	: data1 <= weights[1150];
				12'd1151	: data1 <= weights[1151];
				12'd1152	: data1 <= weights[1152];
				12'd1153	: data1 <= weights[1153];
				12'd1154	: data1 <= weights[1154];
				12'd1155	: data1 <= weights[1155];
				12'd1156	: data1 <= weights[1156];
				12'd1157	: data1 <= weights[1157];
				12'd1158	: data1 <= weights[1158];
				12'd1159	: data1 <= weights[1159];
				12'd1160	: data1 <= weights[1160];
				12'd1161	: data1 <= weights[1161];
				12'd1162	: data1 <= weights[1162];
				12'd1163	: data1 <= weights[1163];
				12'd1164	: data1 <= weights[1164];
				12'd1165	: data1 <= weights[1165];
				12'd1166	: data1 <= weights[1166];
				12'd1167	: data1 <= weights[1167];
				12'd1168	: data1 <= weights[1168];
				12'd1169	: data1 <= weights[1169];
				12'd1170	: data1 <= weights[1170];
				12'd1171	: data1 <= weights[1171];
				12'd1172	: data1 <= weights[1172];
				12'd1173	: data1 <= weights[1173];
				12'd1174	: data1 <= weights[1174];
				12'd1175	: data1 <= weights[1175];
				12'd1176	: data1 <= weights[1176];
				12'd1177	: data1 <= weights[1177];
				12'd1178	: data1 <= weights[1178];
				12'd1179	: data1 <= weights[1179];
				12'd1180	: data1 <= weights[1180];
				12'd1181	: data1 <= weights[1181];
				12'd1182	: data1 <= weights[1182];
				12'd1183	: data1 <= weights[1183];
				12'd1184	: data1 <= weights[1184];
				12'd1185	: data1 <= weights[1185];
				12'd1186	: data1 <= weights[1186];
				12'd1187	: data1 <= weights[1187];
				12'd1188	: data1 <= weights[1188];
				12'd1189	: data1 <= weights[1189];
				12'd1190	: data1 <= weights[1190];
				12'd1191	: data1 <= weights[1191];
				12'd1192	: data1 <= weights[1192];
				12'd1193	: data1 <= weights[1193];
				12'd1194	: data1 <= weights[1194];
				12'd1195	: data1 <= weights[1195];
				12'd1196	: data1 <= weights[1196];
				12'd1197	: data1 <= weights[1197];
				12'd1198	: data1 <= weights[1198];
				12'd1199	: data1 <= weights[1199];
				12'd1200	: data1 <= weights[1200];
				12'd1201	: data1 <= weights[1201];
				12'd1202	: data1 <= weights[1202];
				12'd1203	: data1 <= weights[1203];
				12'd1204	: data1 <= weights[1204];
				12'd1205	: data1 <= weights[1205];
				12'd1206	: data1 <= weights[1206];
				12'd1207	: data1 <= weights[1207];
				12'd1208	: data1 <= weights[1208];
				12'd1209	: data1 <= weights[1209];
				12'd1210	: data1 <= weights[1210];
				12'd1211	: data1 <= weights[1211];
				12'd1212	: data1 <= weights[1212];
				12'd1213	: data1 <= weights[1213];
				12'd1214	: data1 <= weights[1214];
				12'd1215	: data1 <= weights[1215];
				12'd1216	: data1 <= weights[1216];
				12'd1217	: data1 <= weights[1217];
				12'd1218	: data1 <= weights[1218];
				12'd1219	: data1 <= weights[1219];
				12'd1220	: data1 <= weights[1220];
				12'd1221	: data1 <= weights[1221];
				12'd1222	: data1 <= weights[1222];
				12'd1223	: data1 <= weights[1223];
				12'd1224	: data1 <= weights[1224];
				12'd1225	: data1 <= weights[1225];
				12'd1226	: data1 <= weights[1226];
				12'd1227	: data1 <= weights[1227];
				12'd1228	: data1 <= weights[1228];
				12'd1229	: data1 <= weights[1229];
				12'd1230	: data1 <= weights[1230];
				12'd1231	: data1 <= weights[1231];
				12'd1232	: data1 <= weights[1232];
				12'd1233	: data1 <= weights[1233];
				12'd1234	: data1 <= weights[1234];
				12'd1235	: data1 <= weights[1235];
				12'd1236	: data1 <= weights[1236];
				12'd1237	: data1 <= weights[1237];
				12'd1238	: data1 <= weights[1238];
				12'd1239	: data1 <= weights[1239];
				12'd1240	: data1 <= weights[1240];
				12'd1241	: data1 <= weights[1241];
				12'd1242	: data1 <= weights[1242];
				12'd1243	: data1 <= weights[1243];
				12'd1244	: data1 <= weights[1244];
				12'd1245	: data1 <= weights[1245];
				12'd1246	: data1 <= weights[1246];
				12'd1247	: data1 <= weights[1247];
				12'd1248	: data1 <= weights[1248];
				12'd1249	: data1 <= weights[1249];
				12'd1250	: data1 <= weights[1250];
				12'd1251	: data1 <= weights[1251];
				12'd1252	: data1 <= weights[1252];
				12'd1253	: data1 <= weights[1253];
				12'd1254	: data1 <= weights[1254];
				12'd1255	: data1 <= weights[1255];
				12'd1256	: data1 <= weights[1256];
				12'd1257	: data1 <= weights[1257];
				12'd1258	: data1 <= weights[1258];
				12'd1259	: data1 <= weights[1259];
				12'd1260	: data1 <= weights[1260];
				12'd1261	: data1 <= weights[1261];
				12'd1262	: data1 <= weights[1262];
				12'd1263	: data1 <= weights[1263];
				12'd1264	: data1 <= weights[1264];
				12'd1265	: data1 <= weights[1265];
				12'd1266	: data1 <= weights[1266];
				12'd1267	: data1 <= weights[1267];
				12'd1268	: data1 <= weights[1268];
				12'd1269	: data1 <= weights[1269];
				12'd1270	: data1 <= weights[1270];
				12'd1271	: data1 <= weights[1271];
				12'd1272	: data1 <= weights[1272];
				12'd1273	: data1 <= weights[1273];
				12'd1274	: data1 <= weights[1274];
				12'd1275	: data1 <= weights[1275];
				12'd1276	: data1 <= weights[1276];
				12'd1277	: data1 <= weights[1277];
				12'd1278	: data1 <= weights[1278];
				12'd1279	: data1 <= weights[1279];
				12'd1280	: data1 <= weights[1280];
				12'd1281	: data1 <= weights[1281];
				12'd1282	: data1 <= weights[1282];
				12'd1283	: data1 <= weights[1283];
				12'd1284	: data1 <= weights[1284];
				12'd1285	: data1 <= weights[1285];
				12'd1286	: data1 <= weights[1286];
				12'd1287	: data1 <= weights[1287];
				12'd1288	: data1 <= weights[1288];
				12'd1289	: data1 <= weights[1289];
				12'd1290	: data1 <= weights[1290];
				12'd1291	: data1 <= weights[1291];
				12'd1292	: data1 <= weights[1292];
				12'd1293	: data1 <= weights[1293];
				12'd1294	: data1 <= weights[1294];
				12'd1295	: data1 <= weights[1295];
				12'd1296	: data1 <= weights[1296];
				12'd1297	: data1 <= weights[1297];
				12'd1298	: data1 <= weights[1298];
				12'd1299	: data1 <= weights[1299];
				12'd1300	: data1 <= weights[1300];
				12'd1301	: data1 <= weights[1301];
				12'd1302	: data1 <= weights[1302];
				12'd1303	: data1 <= weights[1303];
				12'd1304	: data1 <= weights[1304];
				12'd1305	: data1 <= weights[1305];
				12'd1306	: data1 <= weights[1306];
				12'd1307	: data1 <= weights[1307];
				12'd1308	: data1 <= weights[1308];
				12'd1309	: data1 <= weights[1309];
				12'd1310	: data1 <= weights[1310];
				12'd1311	: data1 <= weights[1311];
				12'd1312	: data1 <= weights[1312];
				12'd1313	: data1 <= weights[1313];
				12'd1314	: data1 <= weights[1314];
				12'd1315	: data1 <= weights[1315];
				12'd1316	: data1 <= weights[1316];
				12'd1317	: data1 <= weights[1317];
				12'd1318	: data1 <= weights[1318];
				12'd1319	: data1 <= weights[1319];
				12'd1320	: data1 <= weights[1320];
				12'd1321	: data1 <= weights[1321];
				12'd1322	: data1 <= weights[1322];
				12'd1323	: data1 <= weights[1323];
				12'd1324	: data1 <= weights[1324];
				12'd1325	: data1 <= weights[1325];
				12'd1326	: data1 <= weights[1326];
				12'd1327	: data1 <= weights[1327];
				12'd1328	: data1 <= weights[1328];
				12'd1329	: data1 <= weights[1329];
				12'd1330	: data1 <= weights[1330];
				12'd1331	: data1 <= weights[1331];
				12'd1332	: data1 <= weights[1332];
				12'd1333	: data1 <= weights[1333];
				12'd1334	: data1 <= weights[1334];
				12'd1335	: data1 <= weights[1335];
				12'd1336	: data1 <= weights[1336];
				12'd1337	: data1 <= weights[1337];
				12'd1338	: data1 <= weights[1338];
				12'd1339	: data1 <= weights[1339];
				12'd1340	: data1 <= weights[1340];
				12'd1341	: data1 <= weights[1341];
				12'd1342	: data1 <= weights[1342];
				12'd1343	: data1 <= weights[1343];
				12'd1344	: data1 <= weights[1344];
				12'd1345	: data1 <= weights[1345];
				12'd1346	: data1 <= weights[1346];
				12'd1347	: data1 <= weights[1347];
				12'd1348	: data1 <= weights[1348];
				12'd1349	: data1 <= weights[1349];
				12'd1350	: data1 <= weights[1350];
				12'd1351	: data1 <= weights[1351];
				12'd1352	: data1 <= weights[1352];
				12'd1353	: data1 <= weights[1353];
				12'd1354	: data1 <= weights[1354];
				12'd1355	: data1 <= weights[1355];
				12'd1356	: data1 <= weights[1356];
				12'd1357	: data1 <= weights[1357];
				12'd1358	: data1 <= weights[1358];
				12'd1359	: data1 <= weights[1359];
				12'd1360	: data1 <= weights[1360];
				12'd1361	: data1 <= weights[1361];
				12'd1362	: data1 <= weights[1362];
				12'd1363	: data1 <= weights[1363];
				12'd1364	: data1 <= weights[1364];
				12'd1365	: data1 <= weights[1365];
				12'd1366	: data1 <= weights[1366];
				12'd1367	: data1 <= weights[1367];
				12'd1368	: data1 <= weights[1368];
				12'd1369	: data1 <= weights[1369];
				12'd1370	: data1 <= weights[1370];
				12'd1371	: data1 <= weights[1371];
				12'd1372	: data1 <= weights[1372];
				12'd1373	: data1 <= weights[1373];
				12'd1374	: data1 <= weights[1374];
				12'd1375	: data1 <= weights[1375];
				12'd1376	: data1 <= weights[1376];
				12'd1377	: data1 <= weights[1377];
				12'd1378	: data1 <= weights[1378];
				12'd1379	: data1 <= weights[1379];
				12'd1380	: data1 <= weights[1380];
				12'd1381	: data1 <= weights[1381];
				12'd1382	: data1 <= weights[1382];
				12'd1383	: data1 <= weights[1383];
				12'd1384	: data1 <= weights[1384];
				12'd1385	: data1 <= weights[1385];
				12'd1386	: data1 <= weights[1386];
				12'd1387	: data1 <= weights[1387];
				12'd1388	: data1 <= weights[1388];
				12'd1389	: data1 <= weights[1389];
				12'd1390	: data1 <= weights[1390];
				12'd1391	: data1 <= weights[1391];
				12'd1392	: data1 <= weights[1392];
				12'd1393	: data1 <= weights[1393];
				12'd1394	: data1 <= weights[1394];
				12'd1395	: data1 <= weights[1395];
				12'd1396	: data1 <= weights[1396];
				12'd1397	: data1 <= weights[1397];
				12'd1398	: data1 <= weights[1398];
				12'd1399	: data1 <= weights[1399];
				12'd1400	: data1 <= weights[1400];
				12'd1401	: data1 <= weights[1401];
				12'd1402	: data1 <= weights[1402];
				12'd1403	: data1 <= weights[1403];
				12'd1404	: data1 <= weights[1404];
				12'd1405	: data1 <= weights[1405];
				12'd1406	: data1 <= weights[1406];
				12'd1407	: data1 <= weights[1407];
				12'd1408	: data1 <= weights[1408];
				12'd1409	: data1 <= weights[1409];
				12'd1410	: data1 <= weights[1410];
				12'd1411	: data1 <= weights[1411];
				12'd1412	: data1 <= weights[1412];
				12'd1413	: data1 <= weights[1413];
				12'd1414	: data1 <= weights[1414];
				12'd1415	: data1 <= weights[1415];
				12'd1416	: data1 <= weights[1416];
				12'd1417	: data1 <= weights[1417];
				12'd1418	: data1 <= weights[1418];
				12'd1419	: data1 <= weights[1419];
				12'd1420	: data1 <= weights[1420];
				12'd1421	: data1 <= weights[1421];
				12'd1422	: data1 <= weights[1422];
				12'd1423	: data1 <= weights[1423];
				12'd1424	: data1 <= weights[1424];
				12'd1425	: data1 <= weights[1425];
				12'd1426	: data1 <= weights[1426];
				12'd1427	: data1 <= weights[1427];
				12'd1428	: data1 <= weights[1428];
				12'd1429	: data1 <= weights[1429];
				12'd1430	: data1 <= weights[1430];
				12'd1431	: data1 <= weights[1431];
				12'd1432	: data1 <= weights[1432];
				12'd1433	: data1 <= weights[1433];
				12'd1434	: data1 <= weights[1434];
				12'd1435	: data1 <= weights[1435];
				12'd1436	: data1 <= weights[1436];
				12'd1437	: data1 <= weights[1437];
				12'd1438	: data1 <= weights[1438];
				12'd1439	: data1 <= weights[1439];
				12'd1440	: data1 <= weights[1440];
				12'd1441	: data1 <= weights[1441];
				12'd1442	: data1 <= weights[1442];
				12'd1443	: data1 <= weights[1443];
				12'd1444	: data1 <= weights[1444];
				12'd1445	: data1 <= weights[1445];
				12'd1446	: data1 <= weights[1446];
				12'd1447	: data1 <= weights[1447];
				12'd1448	: data1 <= weights[1448];
				12'd1449	: data1 <= weights[1449];
				12'd1450	: data1 <= weights[1450];
				12'd1451	: data1 <= weights[1451];
				12'd1452	: data1 <= weights[1452];
				12'd1453	: data1 <= weights[1453];
				12'd1454	: data1 <= weights[1454];
				12'd1455	: data1 <= weights[1455];
				12'd1456	: data1 <= weights[1456];
				12'd1457	: data1 <= weights[1457];
				12'd1458	: data1 <= weights[1458];
				12'd1459	: data1 <= weights[1459];
				12'd1460	: data1 <= weights[1460];
				12'd1461	: data1 <= weights[1461];
				12'd1462	: data1 <= weights[1462];
				12'd1463	: data1 <= weights[1463];
				12'd1464	: data1 <= weights[1464];
				12'd1465	: data1 <= weights[1465];
				12'd1466	: data1 <= weights[1466];
				12'd1467	: data1 <= weights[1467];
				12'd1468	: data1 <= weights[1468];
				12'd1469	: data1 <= weights[1469];
				12'd1470	: data1 <= weights[1470];
				12'd1471	: data1 <= weights[1471];
				12'd1472	: data1 <= weights[1472];
				12'd1473	: data1 <= weights[1473];
				12'd1474	: data1 <= weights[1474];
				12'd1475	: data1 <= weights[1475];
				12'd1476	: data1 <= weights[1476];
				12'd1477	: data1 <= weights[1477];
				12'd1478	: data1 <= weights[1478];
				12'd1479	: data1 <= weights[1479];
				12'd1480	: data1 <= weights[1480];
				12'd1481	: data1 <= weights[1481];
				12'd1482	: data1 <= weights[1482];
				12'd1483	: data1 <= weights[1483];
				12'd1484	: data1 <= weights[1484];
				12'd1485	: data1 <= weights[1485];
				12'd1486	: data1 <= weights[1486];
				12'd1487	: data1 <= weights[1487];
				12'd1488	: data1 <= weights[1488];
				12'd1489	: data1 <= weights[1489];
				12'd1490	: data1 <= weights[1490];
				12'd1491	: data1 <= weights[1491];
				12'd1492	: data1 <= weights[1492];
				12'd1493	: data1 <= weights[1493];
				12'd1494	: data1 <= weights[1494];
				12'd1495	: data1 <= weights[1495];
				12'd1496	: data1 <= weights[1496];
				12'd1497	: data1 <= weights[1497];
				12'd1498	: data1 <= weights[1498];
				12'd1499	: data1 <= weights[1499];
				12'd1500	: data1 <= weights[1500];
				12'd1501	: data1 <= weights[1501];
				12'd1502	: data1 <= weights[1502];
				12'd1503	: data1 <= weights[1503];
				12'd1504	: data1 <= weights[1504];
				12'd1505	: data1 <= weights[1505];
				12'd1506	: data1 <= weights[1506];
				12'd1507	: data1 <= weights[1507];
				12'd1508	: data1 <= weights[1508];
				12'd1509	: data1 <= weights[1509];
				12'd1510	: data1 <= weights[1510];
				12'd1511	: data1 <= weights[1511];
				12'd1512	: data1 <= weights[1512];
				12'd1513	: data1 <= weights[1513];
				12'd1514	: data1 <= weights[1514];
				12'd1515	: data1 <= weights[1515];
				12'd1516	: data1 <= weights[1516];
				12'd1517	: data1 <= weights[1517];
				12'd1518	: data1 <= weights[1518];
				12'd1519	: data1 <= weights[1519];
				12'd1520	: data1 <= weights[1520];
				12'd1521	: data1 <= weights[1521];
				12'd1522	: data1 <= weights[1522];
				12'd1523	: data1 <= weights[1523];
				12'd1524	: data1 <= weights[1524];
				12'd1525	: data1 <= weights[1525];
				12'd1526	: data1 <= weights[1526];
				12'd1527	: data1 <= weights[1527];
				12'd1528	: data1 <= weights[1528];
				12'd1529	: data1 <= weights[1529];
				12'd1530	: data1 <= weights[1530];
				12'd1531	: data1 <= weights[1531];
				12'd1532	: data1 <= weights[1532];
				12'd1533	: data1 <= weights[1533];
				12'd1534	: data1 <= weights[1534];
				12'd1535	: data1 <= weights[1535];
				12'd1536	: data1 <= weights[1536];
				12'd1537	: data1 <= weights[1537];
				12'd1538	: data1 <= weights[1538];
				12'd1539	: data1 <= weights[1539];
				12'd1540	: data1 <= weights[1540];
				12'd1541	: data1 <= weights[1541];
				12'd1542	: data1 <= weights[1542];
				12'd1543	: data1 <= weights[1543];
				12'd1544	: data1 <= weights[1544];
				12'd1545	: data1 <= weights[1545];
				12'd1546	: data1 <= weights[1546];
				12'd1547	: data1 <= weights[1547];
				12'd1548	: data1 <= weights[1548];
				12'd1549	: data1 <= weights[1549];
				12'd1550	: data1 <= weights[1550];
				12'd1551	: data1 <= weights[1551];
				12'd1552	: data1 <= weights[1552];
				12'd1553	: data1 <= weights[1553];
				12'd1554	: data1 <= weights[1554];
				12'd1555	: data1 <= weights[1555];
				12'd1556	: data1 <= weights[1556];
				12'd1557	: data1 <= weights[1557];
				12'd1558	: data1 <= weights[1558];
				12'd1559	: data1 <= weights[1559];
				12'd1560	: data1 <= weights[1560];
				12'd1561	: data1 <= weights[1561];
				12'd1562	: data1 <= weights[1562];
				12'd1563	: data1 <= weights[1563];
				12'd1564	: data1 <= weights[1564];
				12'd1565	: data1 <= weights[1565];
				12'd1566	: data1 <= weights[1566];
				12'd1567	: data1 <= weights[1567];
				12'd1568	: data1 <= weights[1568];
				12'd1569	: data1 <= weights[1569];
				12'd1570	: data1 <= weights[1570];
				12'd1571	: data1 <= weights[1571];
				12'd1572	: data1 <= weights[1572];
				12'd1573	: data1 <= weights[1573];
				12'd1574	: data1 <= weights[1574];
				12'd1575	: data1 <= weights[1575];
				12'd1576	: data1 <= weights[1576];
				12'd1577	: data1 <= weights[1577];
				12'd1578	: data1 <= weights[1578];
				12'd1579	: data1 <= weights[1579];
				12'd1580	: data1 <= weights[1580];
				12'd1581	: data1 <= weights[1581];
				12'd1582	: data1 <= weights[1582];
				12'd1583	: data1 <= weights[1583];
				12'd1584	: data1 <= weights[1584];
				12'd1585	: data1 <= weights[1585];
				12'd1586	: data1 <= weights[1586];
				12'd1587	: data1 <= weights[1587];
				12'd1588	: data1 <= weights[1588];
				12'd1589	: data1 <= weights[1589];
				12'd1590	: data1 <= weights[1590];
				12'd1591	: data1 <= weights[1591];
				12'd1592	: data1 <= weights[1592];
				12'd1593	: data1 <= weights[1593];
				12'd1594	: data1 <= weights[1594];
				12'd1595	: data1 <= weights[1595];
				12'd1596	: data1 <= weights[1596];
				12'd1597	: data1 <= weights[1597];
				12'd1598	: data1 <= weights[1598];
				12'd1599	: data1 <= weights[1599];
				12'd1600	: data1 <= weights[1600];
				12'd1601	: data1 <= weights[1601];
				12'd1602	: data1 <= weights[1602];
				12'd1603	: data1 <= weights[1603];
				12'd1604	: data1 <= weights[1604];
				12'd1605	: data1 <= weights[1605];
				12'd1606	: data1 <= weights[1606];
				12'd1607	: data1 <= weights[1607];
				12'd1608	: data1 <= weights[1608];
				12'd1609	: data1 <= weights[1609];
				12'd1610	: data1 <= weights[1610];
				12'd1611	: data1 <= weights[1611];
				12'd1612	: data1 <= weights[1612];
				12'd1613	: data1 <= weights[1613];
				12'd1614	: data1 <= weights[1614];
				12'd1615	: data1 <= weights[1615];
				12'd1616	: data1 <= weights[1616];
				12'd1617	: data1 <= weights[1617];
				12'd1618	: data1 <= weights[1618];
				12'd1619	: data1 <= weights[1619];
				12'd1620	: data1 <= weights[1620];
				12'd1621	: data1 <= weights[1621];
				12'd1622	: data1 <= weights[1622];
				12'd1623	: data1 <= weights[1623];
				12'd1624	: data1 <= weights[1624];
				12'd1625	: data1 <= weights[1625];
				12'd1626	: data1 <= weights[1626];
				12'd1627	: data1 <= weights[1627];
				12'd1628	: data1 <= weights[1628];
				12'd1629	: data1 <= weights[1629];
				12'd1630	: data1 <= weights[1630];
				12'd1631	: data1 <= weights[1631];
				12'd1632	: data1 <= weights[1632];
				12'd1633	: data1 <= weights[1633];
				12'd1634	: data1 <= weights[1634];
				12'd1635	: data1 <= weights[1635];
				12'd1636	: data1 <= weights[1636];
				12'd1637	: data1 <= weights[1637];
				12'd1638	: data1 <= weights[1638];
				12'd1639	: data1 <= weights[1639];
				12'd1640	: data1 <= weights[1640];
				12'd1641	: data1 <= weights[1641];
				12'd1642	: data1 <= weights[1642];
				12'd1643	: data1 <= weights[1643];
				12'd1644	: data1 <= weights[1644];
				12'd1645	: data1 <= weights[1645];
				12'd1646	: data1 <= weights[1646];
				12'd1647	: data1 <= weights[1647];
				12'd1648	: data1 <= weights[1648];
				12'd1649	: data1 <= weights[1649];
				12'd1650	: data1 <= weights[1650];
				12'd1651	: data1 <= weights[1651];
				12'd1652	: data1 <= weights[1652];
				12'd1653	: data1 <= weights[1653];
				12'd1654	: data1 <= weights[1654];
				12'd1655	: data1 <= weights[1655];
				12'd1656	: data1 <= weights[1656];
				12'd1657	: data1 <= weights[1657];
				12'd1658	: data1 <= weights[1658];
				12'd1659	: data1 <= weights[1659];
				12'd1660	: data1 <= weights[1660];
				12'd1661	: data1 <= weights[1661];
				12'd1662	: data1 <= weights[1662];
				12'd1663	: data1 <= weights[1663];
				12'd1664	: data1 <= weights[1664];
				12'd1665	: data1 <= weights[1665];
				12'd1666	: data1 <= weights[1666];
				12'd1667	: data1 <= weights[1667];
				12'd1668	: data1 <= weights[1668];
				12'd1669	: data1 <= weights[1669];
				12'd1670	: data1 <= weights[1670];
				12'd1671	: data1 <= weights[1671];
				12'd1672	: data1 <= weights[1672];
				12'd1673	: data1 <= weights[1673];
				12'd1674	: data1 <= weights[1674];
				12'd1675	: data1 <= weights[1675];
				12'd1676	: data1 <= weights[1676];
				12'd1677	: data1 <= weights[1677];
				12'd1678	: data1 <= weights[1678];
				12'd1679	: data1 <= weights[1679];
				12'd1680	: data1 <= weights[1680];
				12'd1681	: data1 <= weights[1681];
				12'd1682	: data1 <= weights[1682];
				12'd1683	: data1 <= weights[1683];
				12'd1684	: data1 <= weights[1684];
				12'd1685	: data1 <= weights[1685];
				12'd1686	: data1 <= weights[1686];
				12'd1687	: data1 <= weights[1687];
				12'd1688	: data1 <= weights[1688];
				12'd1689	: data1 <= weights[1689];
				12'd1690	: data1 <= weights[1690];
				12'd1691	: data1 <= weights[1691];
				12'd1692	: data1 <= weights[1692];
				12'd1693	: data1 <= weights[1693];
				12'd1694	: data1 <= weights[1694];
				12'd1695	: data1 <= weights[1695];
				12'd1696	: data1 <= weights[1696];
				12'd1697	: data1 <= weights[1697];
				12'd1698	: data1 <= weights[1698];
				12'd1699	: data1 <= weights[1699];
				12'd1700	: data1 <= weights[1700];
				12'd1701	: data1 <= weights[1701];
				12'd1702	: data1 <= weights[1702];
				12'd1703	: data1 <= weights[1703];
				12'd1704	: data1 <= weights[1704];
				12'd1705	: data1 <= weights[1705];
				12'd1706	: data1 <= weights[1706];
				12'd1707	: data1 <= weights[1707];
				12'd1708	: data1 <= weights[1708];
				12'd1709	: data1 <= weights[1709];
				12'd1710	: data1 <= weights[1710];
				12'd1711	: data1 <= weights[1711];
				12'd1712	: data1 <= weights[1712];
				12'd1713	: data1 <= weights[1713];
				12'd1714	: data1 <= weights[1714];
				12'd1715	: data1 <= weights[1715];
				12'd1716	: data1 <= weights[1716];
				12'd1717	: data1 <= weights[1717];
				12'd1718	: data1 <= weights[1718];
				12'd1719	: data1 <= weights[1719];
				12'd1720	: data1 <= weights[1720];
				12'd1721	: data1 <= weights[1721];
				12'd1722	: data1 <= weights[1722];
				12'd1723	: data1 <= weights[1723];
				12'd1724	: data1 <= weights[1724];
				12'd1725	: data1 <= weights[1725];
				12'd1726	: data1 <= weights[1726];
				12'd1727	: data1 <= weights[1727];
				12'd1728	: data1 <= weights[1728];
				12'd1729	: data1 <= weights[1729];
				12'd1730	: data1 <= weights[1730];
				12'd1731	: data1 <= weights[1731];
				12'd1732	: data1 <= weights[1732];
				12'd1733	: data1 <= weights[1733];
				12'd1734	: data1 <= weights[1734];
				12'd1735	: data1 <= weights[1735];
				12'd1736	: data1 <= weights[1736];
				12'd1737	: data1 <= weights[1737];
				12'd1738	: data1 <= weights[1738];
				12'd1739	: data1 <= weights[1739];
				12'd1740	: data1 <= weights[1740];
				12'd1741	: data1 <= weights[1741];
				12'd1742	: data1 <= weights[1742];
				12'd1743	: data1 <= weights[1743];
				12'd1744	: data1 <= weights[1744];
				12'd1745	: data1 <= weights[1745];
				12'd1746	: data1 <= weights[1746];
				12'd1747	: data1 <= weights[1747];
				12'd1748	: data1 <= weights[1748];
				12'd1749	: data1 <= weights[1749];
				12'd1750	: data1 <= weights[1750];
				12'd1751	: data1 <= weights[1751];
				12'd1752	: data1 <= weights[1752];
				12'd1753	: data1 <= weights[1753];
				12'd1754	: data1 <= weights[1754];
				12'd1755	: data1 <= weights[1755];
				12'd1756	: data1 <= weights[1756];
				12'd1757	: data1 <= weights[1757];
				12'd1758	: data1 <= weights[1758];
				12'd1759	: data1 <= weights[1759];
				12'd1760	: data1 <= weights[1760];
				12'd1761	: data1 <= weights[1761];
				12'd1762	: data1 <= weights[1762];
				12'd1763	: data1 <= weights[1763];
				12'd1764	: data1 <= weights[1764];
				12'd1765	: data1 <= weights[1765];
				12'd1766	: data1 <= weights[1766];
				12'd1767	: data1 <= weights[1767];
				12'd1768	: data1 <= weights[1768];
				12'd1769	: data1 <= weights[1769];
				12'd1770	: data1 <= weights[1770];
				12'd1771	: data1 <= weights[1771];
				12'd1772	: data1 <= weights[1772];
				12'd1773	: data1 <= weights[1773];
				12'd1774	: data1 <= weights[1774];
				12'd1775	: data1 <= weights[1775];
				12'd1776	: data1 <= weights[1776];
				12'd1777	: data1 <= weights[1777];
				12'd1778	: data1 <= weights[1778];
				12'd1779	: data1 <= weights[1779];
				12'd1780	: data1 <= weights[1780];
				12'd1781	: data1 <= weights[1781];
				12'd1782	: data1 <= weights[1782];
				12'd1783	: data1 <= weights[1783];
				12'd1784	: data1 <= weights[1784];
				12'd1785	: data1 <= weights[1785];
				12'd1786	: data1 <= weights[1786];
				12'd1787	: data1 <= weights[1787];
				12'd1788	: data1 <= weights[1788];
				12'd1789	: data1 <= weights[1789];
				12'd1790	: data1 <= weights[1790];
				12'd1791	: data1 <= weights[1791];
				12'd1792	: data1 <= weights[1792];
				12'd1793	: data1 <= weights[1793];
				12'd1794	: data1 <= weights[1794];
				12'd1795	: data1 <= weights[1795];
				12'd1796	: data1 <= weights[1796];
				12'd1797	: data1 <= weights[1797];
				12'd1798	: data1 <= weights[1798];
				12'd1799	: data1 <= weights[1799];
				12'd1800	: data1 <= weights[1800];
				12'd1801	: data1 <= weights[1801];
				12'd1802	: data1 <= weights[1802];
				12'd1803	: data1 <= weights[1803];
				12'd1804	: data1 <= weights[1804];
				12'd1805	: data1 <= weights[1805];
				12'd1806	: data1 <= weights[1806];
				12'd1807	: data1 <= weights[1807];
				12'd1808	: data1 <= weights[1808];
				12'd1809	: data1 <= weights[1809];
				12'd1810	: data1 <= weights[1810];
				12'd1811	: data1 <= weights[1811];
				12'd1812	: data1 <= weights[1812];
				12'd1813	: data1 <= weights[1813];
				12'd1814	: data1 <= weights[1814];
				12'd1815	: data1 <= weights[1815];
				12'd1816	: data1 <= weights[1816];
				12'd1817	: data1 <= weights[1817];
				12'd1818	: data1 <= weights[1818];
				12'd1819	: data1 <= weights[1819];
				12'd1820	: data1 <= weights[1820];
				12'd1821	: data1 <= weights[1821];
				12'd1822	: data1 <= weights[1822];
				12'd1823	: data1 <= weights[1823];
				12'd1824	: data1 <= weights[1824];
				12'd1825	: data1 <= weights[1825];
				12'd1826	: data1 <= weights[1826];
				12'd1827	: data1 <= weights[1827];
				12'd1828	: data1 <= weights[1828];
				12'd1829	: data1 <= weights[1829];
				12'd1830	: data1 <= weights[1830];
				12'd1831	: data1 <= weights[1831];
				12'd1832	: data1 <= weights[1832];
				12'd1833	: data1 <= weights[1833];
				12'd1834	: data1 <= weights[1834];
				12'd1835	: data1 <= weights[1835];
				12'd1836	: data1 <= weights[1836];
				12'd1837	: data1 <= weights[1837];
				12'd1838	: data1 <= weights[1838];
				12'd1839	: data1 <= weights[1839];
				12'd1840	: data1 <= weights[1840];
				12'd1841	: data1 <= weights[1841];
				12'd1842	: data1 <= weights[1842];
				12'd1843	: data1 <= weights[1843];
				12'd1844	: data1 <= weights[1844];
				12'd1845	: data1 <= weights[1845];
				12'd1846	: data1 <= weights[1846];
				12'd1847	: data1 <= weights[1847];
				12'd1848	: data1 <= weights[1848];
				12'd1849	: data1 <= weights[1849];
				12'd1850	: data1 <= weights[1850];
				12'd1851	: data1 <= weights[1851];
				12'd1852	: data1 <= weights[1852];
				12'd1853	: data1 <= weights[1853];
				12'd1854	: data1 <= weights[1854];
				12'd1855	: data1 <= weights[1855];
				12'd1856	: data1 <= weights[1856];
				12'd1857	: data1 <= weights[1857];
				12'd1858	: data1 <= weights[1858];
				12'd1859	: data1 <= weights[1859];
				12'd1860	: data1 <= weights[1860];
				12'd1861	: data1 <= weights[1861];
				12'd1862	: data1 <= weights[1862];
				12'd1863	: data1 <= weights[1863];
				12'd1864	: data1 <= weights[1864];
				12'd1865	: data1 <= weights[1865];
				12'd1866	: data1 <= weights[1866];
				12'd1867	: data1 <= weights[1867];
				12'd1868	: data1 <= weights[1868];
				12'd1869	: data1 <= weights[1869];
				12'd1870	: data1 <= weights[1870];
				12'd1871	: data1 <= weights[1871];
				12'd1872	: data1 <= weights[1872];
				12'd1873	: data1 <= weights[1873];
				12'd1874	: data1 <= weights[1874];
				12'd1875	: data1 <= weights[1875];
				12'd1876	: data1 <= weights[1876];
				12'd1877	: data1 <= weights[1877];
				12'd1878	: data1 <= weights[1878];
				12'd1879	: data1 <= weights[1879];
				12'd1880	: data1 <= weights[1880];
				12'd1881	: data1 <= weights[1881];
				12'd1882	: data1 <= weights[1882];
				12'd1883	: data1 <= weights[1883];
				12'd1884	: data1 <= weights[1884];
				12'd1885	: data1 <= weights[1885];
				12'd1886	: data1 <= weights[1886];
				12'd1887	: data1 <= weights[1887];
				12'd1888	: data1 <= weights[1888];
				12'd1889	: data1 <= weights[1889];
				12'd1890	: data1 <= weights[1890];
				12'd1891	: data1 <= weights[1891];
				12'd1892	: data1 <= weights[1892];
				12'd1893	: data1 <= weights[1893];
				12'd1894	: data1 <= weights[1894];
				12'd1895	: data1 <= weights[1895];
				12'd1896	: data1 <= weights[1896];
				12'd1897	: data1 <= weights[1897];
				12'd1898	: data1 <= weights[1898];
				12'd1899	: data1 <= weights[1899];
				12'd1900	: data1 <= weights[1900];
				12'd1901	: data1 <= weights[1901];
				12'd1902	: data1 <= weights[1902];
				12'd1903	: data1 <= weights[1903];
				12'd1904	: data1 <= weights[1904];
				12'd1905	: data1 <= weights[1905];
				12'd1906	: data1 <= weights[1906];
				12'd1907	: data1 <= weights[1907];
				12'd1908	: data1 <= weights[1908];
				12'd1909	: data1 <= weights[1909];
				12'd1910	: data1 <= weights[1910];
				12'd1911	: data1 <= weights[1911];
				12'd1912	: data1 <= weights[1912];
				12'd1913	: data1 <= weights[1913];
				12'd1914	: data1 <= weights[1914];
				12'd1915	: data1 <= weights[1915];
				12'd1916	: data1 <= weights[1916];
				12'd1917	: data1 <= weights[1917];
				12'd1918	: data1 <= weights[1918];
				12'd1919	: data1 <= weights[1919];
				12'd1920	: data1 <= weights[1920];
				12'd1921	: data1 <= weights[1921];
				12'd1922	: data1 <= weights[1922];
				12'd1923	: data1 <= weights[1923];
				12'd1924	: data1 <= weights[1924];
				12'd1925	: data1 <= weights[1925];
				12'd1926	: data1 <= weights[1926];
				12'd1927	: data1 <= weights[1927];
				12'd1928	: data1 <= weights[1928];
				12'd1929	: data1 <= weights[1929];
				12'd1930	: data1 <= weights[1930];
				12'd1931	: data1 <= weights[1931];
				12'd1932	: data1 <= weights[1932];
				12'd1933	: data1 <= weights[1933];
				12'd1934	: data1 <= weights[1934];
				12'd1935	: data1 <= weights[1935];
				12'd1936	: data1 <= weights[1936];
				12'd1937	: data1 <= weights[1937];
				12'd1938	: data1 <= weights[1938];
				12'd1939	: data1 <= weights[1939];
				12'd1940	: data1 <= weights[1940];
				12'd1941	: data1 <= weights[1941];
				12'd1942	: data1 <= weights[1942];
				12'd1943	: data1 <= weights[1943];
				12'd1944	: data1 <= weights[1944];
				12'd1945	: data1 <= weights[1945];
				12'd1946	: data1 <= weights[1946];
				12'd1947	: data1 <= weights[1947];
				12'd1948	: data1 <= weights[1948];
				12'd1949	: data1 <= weights[1949];
				12'd1950	: data1 <= weights[1950];
				12'd1951	: data1 <= weights[1951];
				12'd1952	: data1 <= weights[1952];
				12'd1953	: data1 <= weights[1953];
				12'd1954	: data1 <= weights[1954];
				12'd1955	: data1 <= weights[1955];
				12'd1956	: data1 <= weights[1956];
				12'd1957	: data1 <= weights[1957];
				12'd1958	: data1 <= weights[1958];
				12'd1959	: data1 <= weights[1959];
				12'd1960	: data1 <= weights[1960];
				12'd1961	: data1 <= weights[1961];
				12'd1962	: data1 <= weights[1962];
				12'd1963	: data1 <= weights[1963];
				12'd1964	: data1 <= weights[1964];
				12'd1965	: data1 <= weights[1965];
				12'd1966	: data1 <= weights[1966];
				12'd1967	: data1 <= weights[1967];
				12'd1968	: data1 <= weights[1968];
				12'd1969	: data1 <= weights[1969];
				12'd1970	: data1 <= weights[1970];
				12'd1971	: data1 <= weights[1971];
				12'd1972	: data1 <= weights[1972];
				12'd1973	: data1 <= weights[1973];
				12'd1974	: data1 <= weights[1974];
				12'd1975	: data1 <= weights[1975];
				12'd1976	: data1 <= weights[1976];
				12'd1977	: data1 <= weights[1977];
				12'd1978	: data1 <= weights[1978];
				12'd1979	: data1 <= weights[1979];
				12'd1980	: data1 <= weights[1980];
				12'd1981	: data1 <= weights[1981];
				12'd1982	: data1 <= weights[1982];
				12'd1983	: data1 <= weights[1983];
				12'd1984	: data1 <= weights[1984];
				12'd1985	: data1 <= weights[1985];
				12'd1986	: data1 <= weights[1986];
				12'd1987	: data1 <= weights[1987];
				12'd1988	: data1 <= weights[1988];
				12'd1989	: data1 <= weights[1989];
				12'd1990	: data1 <= weights[1990];
				12'd1991	: data1 <= weights[1991];
				12'd1992	: data1 <= weights[1992];
				12'd1993	: data1 <= weights[1993];
				12'd1994	: data1 <= weights[1994];
				12'd1995	: data1 <= weights[1995];
				12'd1996	: data1 <= weights[1996];
				12'd1997	: data1 <= weights[1997];
				12'd1998	: data1 <= weights[1998];
				12'd1999	: data1 <= weights[1999];
				12'd2000	: data1 <= weights[2000];
				12'd2001	: data1 <= weights[2001];
				12'd2002	: data1 <= weights[2002];
				12'd2003	: data1 <= weights[2003];
				12'd2004	: data1 <= weights[2004];
				12'd2005	: data1 <= weights[2005];
				12'd2006	: data1 <= weights[2006];
				12'd2007	: data1 <= weights[2007];
				12'd2008	: data1 <= weights[2008];
				12'd2009	: data1 <= weights[2009];
				12'd2010	: data1 <= weights[2010];
				12'd2011	: data1 <= weights[2011];
				12'd2012	: data1 <= weights[2012];
				12'd2013	: data1 <= weights[2013];
				12'd2014	: data1 <= weights[2014];
				12'd2015	: data1 <= weights[2015];
				12'd2016	: data1 <= weights[2016];
				12'd2017	: data1 <= weights[2017];
				12'd2018	: data1 <= weights[2018];
				12'd2019	: data1 <= weights[2019];
				12'd2020	: data1 <= weights[2020];
				12'd2021	: data1 <= weights[2021];
				12'd2022	: data1 <= weights[2022];
				12'd2023	: data1 <= weights[2023];
				12'd2024	: data1 <= weights[2024];
				12'd2025	: data1 <= weights[2025];
				12'd2026	: data1 <= weights[2026];
				12'd2027	: data1 <= weights[2027];
				12'd2028	: data1 <= weights[2028];
				12'd2029	: data1 <= weights[2029];
				12'd2030	: data1 <= weights[2030];
				12'd2031	: data1 <= weights[2031];
				12'd2032	: data1 <= weights[2032];
				12'd2033	: data1 <= weights[2033];
				12'd2034	: data1 <= weights[2034];
				12'd2035	: data1 <= weights[2035];
				12'd2036	: data1 <= weights[2036];
				12'd2037	: data1 <= weights[2037];
				12'd2038	: data1 <= weights[2038];
				12'd2039	: data1 <= weights[2039];
				12'd2040	: data1 <= weights[2040];
				12'd2041	: data1 <= weights[2041];
				12'd2042	: data1 <= weights[2042];
				12'd2043	: data1 <= weights[2043];
				12'd2044	: data1 <= weights[2044];
				12'd2045	: data1 <= weights[2045];
				12'd2046	: data1 <= weights[2046];
				12'd2047	: data1 <= weights[2047];
				12'd2048	: data1 <= weights[2048];
				12'd2049	: data1 <= weights[2049];
				12'd2050	: data1 <= weights[2050];
				12'd2051	: data1 <= weights[2051];
				12'd2052	: data1 <= weights[2052];
				12'd2053	: data1 <= weights[2053];
				12'd2054	: data1 <= weights[2054];
				12'd2055	: data1 <= weights[2055];
				12'd2056	: data1 <= weights[2056];
				12'd2057	: data1 <= weights[2057];
				12'd2058	: data1 <= weights[2058];
				12'd2059	: data1 <= weights[2059];
				12'd2060	: data1 <= weights[2060];
				12'd2061	: data1 <= weights[2061];
				12'd2062	: data1 <= weights[2062];
				12'd2063	: data1 <= weights[2063];
				12'd2064	: data1 <= weights[2064];
				12'd2065	: data1 <= weights[2065];
				12'd2066	: data1 <= weights[2066];
				12'd2067	: data1 <= weights[2067];
				12'd2068	: data1 <= weights[2068];
				12'd2069	: data1 <= weights[2069];
				12'd2070	: data1 <= weights[2070];
				12'd2071	: data1 <= weights[2071];
				12'd2072	: data1 <= weights[2072];
				12'd2073	: data1 <= weights[2073];
				12'd2074	: data1 <= weights[2074];
				12'd2075	: data1 <= weights[2075];
				12'd2076	: data1 <= weights[2076];
				12'd2077	: data1 <= weights[2077];
				12'd2078	: data1 <= weights[2078];
				12'd2079	: data1 <= weights[2079];
				12'd2080	: data1 <= weights[2080];
				12'd2081	: data1 <= weights[2081];
				12'd2082	: data1 <= weights[2082];
				12'd2083	: data1 <= weights[2083];
				12'd2084	: data1 <= weights[2084];
				12'd2085	: data1 <= weights[2085];
				12'd2086	: data1 <= weights[2086];
				12'd2087	: data1 <= weights[2087];
				12'd2088	: data1 <= weights[2088];
				12'd2089	: data1 <= weights[2089];
				12'd2090	: data1 <= weights[2090];
				12'd2091	: data1 <= weights[2091];
				12'd2092	: data1 <= weights[2092];
				12'd2093	: data1 <= weights[2093];
				12'd2094	: data1 <= weights[2094];
				12'd2095	: data1 <= weights[2095];
				12'd2096	: data1 <= weights[2096];
				12'd2097	: data1 <= weights[2097];
				12'd2098	: data1 <= weights[2098];
				12'd2099	: data1 <= weights[2099];
				12'd2100	: data1 <= weights[2100];
				12'd2101	: data1 <= weights[2101];
				12'd2102	: data1 <= weights[2102];
				12'd2103	: data1 <= weights[2103];
				12'd2104	: data1 <= weights[2104];
				12'd2105	: data1 <= weights[2105];
				12'd2106	: data1 <= weights[2106];
				12'd2107	: data1 <= weights[2107];
				12'd2108	: data1 <= weights[2108];
				12'd2109	: data1 <= weights[2109];
				12'd2110	: data1 <= weights[2110];
				12'd2111	: data1 <= weights[2111];
				12'd2112	: data1 <= weights[2112];
				12'd2113	: data1 <= weights[2113];
				12'd2114	: data1 <= weights[2114];
				12'd2115	: data1 <= weights[2115];
				12'd2116	: data1 <= weights[2116];
				12'd2117	: data1 <= weights[2117];
				12'd2118	: data1 <= weights[2118];
				12'd2119	: data1 <= weights[2119];
				12'd2120	: data1 <= weights[2120];
				12'd2121	: data1 <= weights[2121];
				12'd2122	: data1 <= weights[2122];
				12'd2123	: data1 <= weights[2123];
				12'd2124	: data1 <= weights[2124];
				12'd2125	: data1 <= weights[2125];
				12'd2126	: data1 <= weights[2126];
				12'd2127	: data1 <= weights[2127];
				12'd2128	: data1 <= weights[2128];
				12'd2129	: data1 <= weights[2129];
				12'd2130	: data1 <= weights[2130];
				12'd2131	: data1 <= weights[2131];
				12'd2132	: data1 <= weights[2132];
				12'd2133	: data1 <= weights[2133];
				12'd2134	: data1 <= weights[2134];
				12'd2135	: data1 <= weights[2135];
				12'd2136	: data1 <= weights[2136];
				12'd2137	: data1 <= weights[2137];
				12'd2138	: data1 <= weights[2138];
				12'd2139	: data1 <= weights[2139];
				12'd2140	: data1 <= weights[2140];
				12'd2141	: data1 <= weights[2141];
				12'd2142	: data1 <= weights[2142];
				12'd2143	: data1 <= weights[2143];
				12'd2144	: data1 <= weights[2144];
				12'd2145	: data1 <= weights[2145];
				12'd2146	: data1 <= weights[2146];
				12'd2147	: data1 <= weights[2147];
				12'd2148	: data1 <= weights[2148];
				12'd2149	: data1 <= weights[2149];
				12'd2150	: data1 <= weights[2150];
				12'd2151	: data1 <= weights[2151];
				12'd2152	: data1 <= weights[2152];
				12'd2153	: data1 <= weights[2153];
				12'd2154	: data1 <= weights[2154];
				12'd2155	: data1 <= weights[2155];
				12'd2156	: data1 <= weights[2156];
				12'd2157	: data1 <= weights[2157];
				12'd2158	: data1 <= weights[2158];
				12'd2159	: data1 <= weights[2159];
				12'd2160	: data1 <= weights[2160];
				12'd2161	: data1 <= weights[2161];
				12'd2162	: data1 <= weights[2162];
				12'd2163	: data1 <= weights[2163];
				12'd2164	: data1 <= weights[2164];
				12'd2165	: data1 <= weights[2165];
				12'd2166	: data1 <= weights[2166];
				12'd2167	: data1 <= weights[2167];
				12'd2168	: data1 <= weights[2168];
				12'd2169	: data1 <= weights[2169];
				12'd2170	: data1 <= weights[2170];
				12'd2171	: data1 <= weights[2171];
				12'd2172	: data1 <= weights[2172];
				12'd2173	: data1 <= weights[2173];
				12'd2174	: data1 <= weights[2174];
				12'd2175	: data1 <= weights[2175];
				12'd2176	: data1 <= weights[2176];
				12'd2177	: data1 <= weights[2177];
				12'd2178	: data1 <= weights[2178];
				12'd2179	: data1 <= weights[2179];
				12'd2180	: data1 <= weights[2180];
				12'd2181	: data1 <= weights[2181];
				12'd2182	: data1 <= weights[2182];
				12'd2183	: data1 <= weights[2183];
				12'd2184	: data1 <= weights[2184];
				12'd2185	: data1 <= weights[2185];
				12'd2186	: data1 <= weights[2186];
				12'd2187	: data1 <= weights[2187];
				12'd2188	: data1 <= weights[2188];
				12'd2189	: data1 <= weights[2189];
				12'd2190	: data1 <= weights[2190];
				12'd2191	: data1 <= weights[2191];
				12'd2192	: data1 <= weights[2192];
				12'd2193	: data1 <= weights[2193];
				12'd2194	: data1 <= weights[2194];
				12'd2195	: data1 <= weights[2195];
				12'd2196	: data1 <= weights[2196];
				12'd2197	: data1 <= weights[2197];
				12'd2198	: data1 <= weights[2198];
				12'd2199	: data1 <= weights[2199];
				12'd2200	: data1 <= weights[2200];
				12'd2201	: data1 <= weights[2201];
				12'd2202	: data1 <= weights[2202];
				12'd2203	: data1 <= weights[2203];
				12'd2204	: data1 <= weights[2204];
				12'd2205	: data1 <= weights[2205];
				12'd2206	: data1 <= weights[2206];
				12'd2207	: data1 <= weights[2207];
				12'd2208	: data1 <= weights[2208];
				12'd2209	: data1 <= weights[2209];
				12'd2210	: data1 <= weights[2210];
				12'd2211	: data1 <= weights[2211];
				12'd2212	: data1 <= weights[2212];
				12'd2213	: data1 <= weights[2213];
				12'd2214	: data1 <= weights[2214];
				12'd2215	: data1 <= weights[2215];
				12'd2216	: data1 <= weights[2216];
				12'd2217	: data1 <= weights[2217];
				12'd2218	: data1 <= weights[2218];
				12'd2219	: data1 <= weights[2219];
				12'd2220	: data1 <= weights[2220];
				12'd2221	: data1 <= weights[2221];
				12'd2222	: data1 <= weights[2222];
				12'd2223	: data1 <= weights[2223];
				12'd2224	: data1 <= weights[2224];
				12'd2225	: data1 <= weights[2225];
				12'd2226	: data1 <= weights[2226];
				12'd2227	: data1 <= weights[2227];
				12'd2228	: data1 <= weights[2228];
				12'd2229	: data1 <= weights[2229];
				12'd2230	: data1 <= weights[2230];
				12'd2231	: data1 <= weights[2231];
				12'd2232	: data1 <= weights[2232];
				12'd2233	: data1 <= weights[2233];
				12'd2234	: data1 <= weights[2234];
				12'd2235	: data1 <= weights[2235];
				12'd2236	: data1 <= weights[2236];
				12'd2237	: data1 <= weights[2237];
				12'd2238	: data1 <= weights[2238];
				12'd2239	: data1 <= weights[2239];
				12'd2240	: data1 <= weights[2240];
				12'd2241	: data1 <= weights[2241];
				12'd2242	: data1 <= weights[2242];
				12'd2243	: data1 <= weights[2243];
				12'd2244	: data1 <= weights[2244];
				12'd2245	: data1 <= weights[2245];
				12'd2246	: data1 <= weights[2246];
				12'd2247	: data1 <= weights[2247];
				12'd2248	: data1 <= weights[2248];
				12'd2249	: data1 <= weights[2249];
				12'd2250	: data1 <= weights[2250];
				12'd2251	: data1 <= weights[2251];
				12'd2252	: data1 <= weights[2252];
				12'd2253	: data1 <= weights[2253];
				12'd2254	: data1 <= weights[2254];
				12'd2255	: data1 <= weights[2255];
				12'd2256	: data1 <= weights[2256];
				12'd2257	: data1 <= weights[2257];
				12'd2258	: data1 <= weights[2258];
				12'd2259	: data1 <= weights[2259];
				12'd2260	: data1 <= weights[2260];
				12'd2261	: data1 <= weights[2261];
				12'd2262	: data1 <= weights[2262];
				12'd2263	: data1 <= weights[2263];
				12'd2264	: data1 <= weights[2264];
				12'd2265	: data1 <= weights[2265];
				12'd2266	: data1 <= weights[2266];
				12'd2267	: data1 <= weights[2267];
				12'd2268	: data1 <= weights[2268];
				12'd2269	: data1 <= weights[2269];
				12'd2270	: data1 <= weights[2270];
				12'd2271	: data1 <= weights[2271];
				12'd2272	: data1 <= weights[2272];
				12'd2273	: data1 <= weights[2273];
				12'd2274	: data1 <= weights[2274];
				12'd2275	: data1 <= weights[2275];
				12'd2276	: data1 <= weights[2276];
				12'd2277	: data1 <= weights[2277];
				12'd2278	: data1 <= weights[2278];
				12'd2279	: data1 <= weights[2279];
				12'd2280	: data1 <= weights[2280];
				12'd2281	: data1 <= weights[2281];
				12'd2282	: data1 <= weights[2282];
				12'd2283	: data1 <= weights[2283];
				12'd2284	: data1 <= weights[2284];
				12'd2285	: data1 <= weights[2285];
				12'd2286	: data1 <= weights[2286];
				12'd2287	: data1 <= weights[2287];
				12'd2288	: data1 <= weights[2288];
				12'd2289	: data1 <= weights[2289];
				12'd2290	: data1 <= weights[2290];
				12'd2291	: data1 <= weights[2291];
				12'd2292	: data1 <= weights[2292];
				12'd2293	: data1 <= weights[2293];
				12'd2294	: data1 <= weights[2294];
				12'd2295	: data1 <= weights[2295];
				12'd2296	: data1 <= weights[2296];
				12'd2297	: data1 <= weights[2297];
				12'd2298	: data1 <= weights[2298];
				12'd2299	: data1 <= weights[2299];
				12'd2300	: data1 <= weights[2300];
				12'd2301	: data1 <= weights[2301];
				12'd2302	: data1 <= weights[2302];
				12'd2303	: data1 <= weights[2303];
				12'd2304	: data1 <= weights[2304];
				12'd2305	: data1 <= weights[2305];
				12'd2306	: data1 <= weights[2306];
				12'd2307	: data1 <= weights[2307];
				12'd2308	: data1 <= weights[2308];
				12'd2309	: data1 <= weights[2309];
				12'd2310	: data1 <= weights[2310];
				12'd2311	: data1 <= weights[2311];
				12'd2312	: data1 <= weights[2312];
				12'd2313	: data1 <= weights[2313];
				12'd2314	: data1 <= weights[2314];
				12'd2315	: data1 <= weights[2315];
				12'd2316	: data1 <= weights[2316];
				12'd2317	: data1 <= weights[2317];
				12'd2318	: data1 <= weights[2318];
				12'd2319	: data1 <= weights[2319];
				12'd2320	: data1 <= weights[2320];
				12'd2321	: data1 <= weights[2321];
				12'd2322	: data1 <= weights[2322];
				12'd2323	: data1 <= weights[2323];
				12'd2324	: data1 <= weights[2324];
				12'd2325	: data1 <= weights[2325];
				12'd2326	: data1 <= weights[2326];
				12'd2327	: data1 <= weights[2327];
				12'd2328	: data1 <= weights[2328];
				12'd2329	: data1 <= weights[2329];
				12'd2330	: data1 <= weights[2330];
				12'd2331	: data1 <= weights[2331];
				12'd2332	: data1 <= weights[2332];
				12'd2333	: data1 <= weights[2333];
				12'd2334	: data1 <= weights[2334];
				12'd2335	: data1 <= weights[2335];
				12'd2336	: data1 <= weights[2336];
				12'd2337	: data1 <= weights[2337];
				12'd2338	: data1 <= weights[2338];
				12'd2339	: data1 <= weights[2339];
				12'd2340	: data1 <= weights[2340];
				12'd2341	: data1 <= weights[2341];
				12'd2342	: data1 <= weights[2342];
				12'd2343	: data1 <= weights[2343];
				12'd2344	: data1 <= weights[2344];
				12'd2345	: data1 <= weights[2345];
				12'd2346	: data1 <= weights[2346];
				12'd2347	: data1 <= weights[2347];
				12'd2348	: data1 <= weights[2348];
				12'd2349	: data1 <= weights[2349];
				12'd2350	: data1 <= weights[2350];
				12'd2351	: data1 <= weights[2351];
				12'd2352	: data1 <= weights[2352];
				12'd2353	: data1 <= weights[2353];
				12'd2354	: data1 <= weights[2354];
				12'd2355	: data1 <= weights[2355];
				12'd2356	: data1 <= weights[2356];
				12'd2357	: data1 <= weights[2357];
				12'd2358	: data1 <= weights[2358];
				12'd2359	: data1 <= weights[2359];
				12'd2360	: data1 <= weights[2360];
				12'd2361	: data1 <= weights[2361];
				12'd2362	: data1 <= weights[2362];
				12'd2363	: data1 <= weights[2363];
				12'd2364	: data1 <= weights[2364];
				12'd2365	: data1 <= weights[2365];
				12'd2366	: data1 <= weights[2366];
				12'd2367	: data1 <= weights[2367];
				12'd2368	: data1 <= weights[2368];
				12'd2369	: data1 <= weights[2369];
				12'd2370	: data1 <= weights[2370];
				12'd2371	: data1 <= weights[2371];
				12'd2372	: data1 <= weights[2372];
				12'd2373	: data1 <= weights[2373];
				12'd2374	: data1 <= weights[2374];
				12'd2375	: data1 <= weights[2375];
				12'd2376	: data1 <= weights[2376];
				12'd2377	: data1 <= weights[2377];
				12'd2378	: data1 <= weights[2378];
				12'd2379	: data1 <= weights[2379];
				12'd2380	: data1 <= weights[2380];
				12'd2381	: data1 <= weights[2381];
				12'd2382	: data1 <= weights[2382];
				12'd2383	: data1 <= weights[2383];
				12'd2384	: data1 <= weights[2384];
				12'd2385	: data1 <= weights[2385];
				12'd2386	: data1 <= weights[2386];
				12'd2387	: data1 <= weights[2387];
				12'd2388	: data1 <= weights[2388];
				12'd2389	: data1 <= weights[2389];
				12'd2390	: data1 <= weights[2390];
				12'd2391	: data1 <= weights[2391];
				12'd2392	: data1 <= weights[2392];
				12'd2393	: data1 <= weights[2393];
				12'd2394	: data1 <= weights[2394];
				12'd2395	: data1 <= weights[2395];
				12'd2396	: data1 <= weights[2396];
				12'd2397	: data1 <= weights[2397];
				12'd2398	: data1 <= weights[2398];
				12'd2399	: data1 <= weights[2399];
				12'd2400	: data1 <= weights[2400];
				12'd2401	: data1 <= weights[2401];
				12'd2402	: data1 <= weights[2402];
				12'd2403	: data1 <= weights[2403];
				12'd2404	: data1 <= weights[2404];
				12'd2405	: data1 <= weights[2405];
				12'd2406	: data1 <= weights[2406];
				12'd2407	: data1 <= weights[2407];
				12'd2408	: data1 <= weights[2408];
				12'd2409	: data1 <= weights[2409];
				12'd2410	: data1 <= weights[2410];
				12'd2411	: data1 <= weights[2411];
				12'd2412	: data1 <= weights[2412];
				12'd2413	: data1 <= weights[2413];
				12'd2414	: data1 <= weights[2414];
				12'd2415	: data1 <= weights[2415];
				12'd2416	: data1 <= weights[2416];
				12'd2417	: data1 <= weights[2417];
				12'd2418	: data1 <= weights[2418];
				12'd2419	: data1 <= weights[2419];
				12'd2420	: data1 <= weights[2420];
				12'd2421	: data1 <= weights[2421];
				12'd2422	: data1 <= weights[2422];
				12'd2423	: data1 <= weights[2423];
				12'd2424	: data1 <= weights[2424];
				12'd2425	: data1 <= weights[2425];
				12'd2426	: data1 <= weights[2426];
				12'd2427	: data1 <= weights[2427];
				12'd2428	: data1 <= weights[2428];
				12'd2429	: data1 <= weights[2429];
				12'd2430	: data1 <= weights[2430];
				12'd2431	: data1 <= weights[2431];
				12'd2432	: data1 <= weights[2432];
				12'd2433	: data1 <= weights[2433];
				12'd2434	: data1 <= weights[2434];
				12'd2435	: data1 <= weights[2435];
				12'd2436	: data1 <= weights[2436];
				12'd2437	: data1 <= weights[2437];
				12'd2438	: data1 <= weights[2438];
				12'd2439	: data1 <= weights[2439];
				12'd2440	: data1 <= weights[2440];
				12'd2441	: data1 <= weights[2441];
				12'd2442	: data1 <= weights[2442];
				12'd2443	: data1 <= weights[2443];
				12'd2444	: data1 <= weights[2444];
				12'd2445	: data1 <= weights[2445];
				12'd2446	: data1 <= weights[2446];
				12'd2447	: data1 <= weights[2447];
				12'd2448	: data1 <= weights[2448];
				12'd2449	: data1 <= weights[2449];
				12'd2450	: data1 <= weights[2450];
				12'd2451	: data1 <= weights[2451];
				12'd2452	: data1 <= weights[2452];
				12'd2453	: data1 <= weights[2453];
				12'd2454	: data1 <= weights[2454];
				12'd2455	: data1 <= weights[2455];
				12'd2456	: data1 <= weights[2456];
				12'd2457	: data1 <= weights[2457];
				12'd2458	: data1 <= weights[2458];
				12'd2459	: data1 <= weights[2459];
				12'd2460	: data1 <= weights[2460];
				12'd2461	: data1 <= weights[2461];
				12'd2462	: data1 <= weights[2462];
				12'd2463	: data1 <= weights[2463];
				12'd2464	: data1 <= weights[2464];
				12'd2465	: data1 <= weights[2465];
				12'd2466	: data1 <= weights[2466];
				12'd2467	: data1 <= weights[2467];
				12'd2468	: data1 <= weights[2468];
				12'd2469	: data1 <= weights[2469];
				12'd2470	: data1 <= weights[2470];
				12'd2471	: data1 <= weights[2471];
				12'd2472	: data1 <= weights[2472];
				12'd2473	: data1 <= weights[2473];
				12'd2474	: data1 <= weights[2474];
				12'd2475	: data1 <= weights[2475];
				12'd2476	: data1 <= weights[2476];
				12'd2477	: data1 <= weights[2477];
				12'd2478	: data1 <= weights[2478];
				12'd2479	: data1 <= weights[2479];
				12'd2480	: data1 <= weights[2480];
				12'd2481	: data1 <= weights[2481];
				12'd2482	: data1 <= weights[2482];
				12'd2483	: data1 <= weights[2483];
				12'd2484	: data1 <= weights[2484];
				12'd2485	: data1 <= weights[2485];
				12'd2486	: data1 <= weights[2486];
				12'd2487	: data1 <= weights[2487];
				12'd2488	: data1 <= weights[2488];
				12'd2489	: data1 <= weights[2489];
				12'd2490	: data1 <= weights[2490];
				12'd2491	: data1 <= weights[2491];
				12'd2492	: data1 <= weights[2492];
				12'd2493	: data1 <= weights[2493];
				12'd2494	: data1 <= weights[2494];
				12'd2495	: data1 <= weights[2495];
				12'd2496	: data1 <= weights[2496];
				12'd2497	: data1 <= weights[2497];
				12'd2498	: data1 <= weights[2498];
				12'd2499	: data1 <= weights[2499];
				12'd2500	: data1 <= weights[2500];
				12'd2501	: data1 <= weights[2501];
				12'd2502	: data1 <= weights[2502];
				12'd2503	: data1 <= weights[2503];
				12'd2504	: data1 <= weights[2504];
				12'd2505	: data1 <= weights[2505];
				12'd2506	: data1 <= weights[2506];
				12'd2507	: data1 <= weights[2507];
				12'd2508	: data1 <= weights[2508];
				12'd2509	: data1 <= weights[2509];
				12'd2510	: data1 <= weights[2510];
				12'd2511	: data1 <= weights[2511];
				12'd2512	: data1 <= weights[2512];
				12'd2513	: data1 <= weights[2513];
				12'd2514	: data1 <= weights[2514];
				12'd2515	: data1 <= weights[2515];
				12'd2516	: data1 <= weights[2516];
				12'd2517	: data1 <= weights[2517];
				12'd2518	: data1 <= weights[2518];
				12'd2519	: data1 <= weights[2519];
				12'd2520	: data1 <= weights[2520];
				12'd2521	: data1 <= weights[2521];
				12'd2522	: data1 <= weights[2522];
				12'd2523	: data1 <= weights[2523];
				12'd2524	: data1 <= weights[2524];
				12'd2525	: data1 <= weights[2525];
				12'd2526	: data1 <= weights[2526];
				12'd2527	: data1 <= weights[2527];
				12'd2528	: data1 <= weights[2528];
				12'd2529	: data1 <= weights[2529];
				12'd2530	: data1 <= weights[2530];
				12'd2531	: data1 <= weights[2531];
				12'd2532	: data1 <= weights[2532];
				12'd2533	: data1 <= weights[2533];
				12'd2534	: data1 <= weights[2534];
				12'd2535	: data1 <= weights[2535];
				12'd2536	: data1 <= weights[2536];
				12'd2537	: data1 <= weights[2537];
				12'd2538	: data1 <= weights[2538];
				12'd2539	: data1 <= weights[2539];
				12'd2540	: data1 <= weights[2540];
				12'd2541	: data1 <= weights[2541];
				12'd2542	: data1 <= weights[2542];
				12'd2543	: data1 <= weights[2543];
				12'd2544	: data1 <= weights[2544];
				12'd2545	: data1 <= weights[2545];
				12'd2546	: data1 <= weights[2546];
				12'd2547	: data1 <= weights[2547];
				12'd2548	: data1 <= weights[2548];
				12'd2549	: data1 <= weights[2549];
				12'd2550	: data1 <= weights[2550];
				12'd2551	: data1 <= weights[2551];
				12'd2552	: data1 <= weights[2552];
				12'd2553	: data1 <= weights[2553];
				12'd2554	: data1 <= weights[2554];
				12'd2555	: data1 <= weights[2555];
				12'd2556	: data1 <= weights[2556];
				12'd2557	: data1 <= weights[2557];
				12'd2558	: data1 <= weights[2558];
				12'd2559	: data1 <= weights[2559];
				12'd2560	: data1 <= weights[2560];
				12'd2561	: data1 <= weights[2561];
				12'd2562	: data1 <= weights[2562];
				12'd2563	: data1 <= weights[2563];
				12'd2564	: data1 <= weights[2564];
				12'd2565	: data1 <= weights[2565];
				12'd2566	: data1 <= weights[2566];
				12'd2567	: data1 <= weights[2567];
				12'd2568	: data1 <= weights[2568];
				12'd2569	: data1 <= weights[2569];
				12'd2570	: data1 <= weights[2570];
				12'd2571	: data1 <= weights[2571];
				12'd2572	: data1 <= weights[2572];
				12'd2573	: data1 <= weights[2573];
				12'd2574	: data1 <= weights[2574];
				12'd2575	: data1 <= weights[2575];
				12'd2576	: data1 <= weights[2576];
				12'd2577	: data1 <= weights[2577];
				12'd2578	: data1 <= weights[2578];
				12'd2579	: data1 <= weights[2579];
				12'd2580	: data1 <= weights[2580];
				12'd2581	: data1 <= weights[2581];
				12'd2582	: data1 <= weights[2582];
				12'd2583	: data1 <= weights[2583];
				12'd2584	: data1 <= weights[2584];
				12'd2585	: data1 <= weights[2585];
				12'd2586	: data1 <= weights[2586];
				12'd2587	: data1 <= weights[2587];
				12'd2588	: data1 <= weights[2588];
				12'd2589	: data1 <= weights[2589];
				12'd2590	: data1 <= weights[2590];
				12'd2591	: data1 <= weights[2591];
				12'd2592	: data1 <= weights[2592];
				12'd2593	: data1 <= weights[2593];
				12'd2594	: data1 <= weights[2594];
				12'd2595	: data1 <= weights[2595];
				12'd2596	: data1 <= weights[2596];
				12'd2597	: data1 <= weights[2597];
				12'd2598	: data1 <= weights[2598];
				12'd2599	: data1 <= weights[2599];
				12'd2600	: data1 <= weights[2600];
				12'd2601	: data1 <= weights[2601];
				12'd2602	: data1 <= weights[2602];
				12'd2603	: data1 <= weights[2603];
				12'd2604	: data1 <= weights[2604];
				12'd2605	: data1 <= weights[2605];
				12'd2606	: data1 <= weights[2606];
				12'd2607	: data1 <= weights[2607];
				12'd2608	: data1 <= weights[2608];
				12'd2609	: data1 <= weights[2609];
				12'd2610	: data1 <= weights[2610];
				12'd2611	: data1 <= weights[2611];
				12'd2612	: data1 <= weights[2612];
				12'd2613	: data1 <= weights[2613];
				12'd2614	: data1 <= weights[2614];
				12'd2615	: data1 <= weights[2615];
				12'd2616	: data1 <= weights[2616];
				12'd2617	: data1 <= weights[2617];
				12'd2618	: data1 <= weights[2618];
				12'd2619	: data1 <= weights[2619];
				12'd2620	: data1 <= weights[2620];
				12'd2621	: data1 <= weights[2621];
				12'd2622	: data1 <= weights[2622];
				12'd2623	: data1 <= weights[2623];
				12'd2624	: data1 <= weights[2624];
				12'd2625	: data1 <= weights[2625];
				12'd2626	: data1 <= weights[2626];
				12'd2627	: data1 <= weights[2627];
				12'd2628	: data1 <= weights[2628];
				12'd2629	: data1 <= weights[2629];
				12'd2630	: data1 <= weights[2630];
				12'd2631	: data1 <= weights[2631];
				12'd2632	: data1 <= weights[2632];
				12'd2633	: data1 <= weights[2633];
				12'd2634	: data1 <= weights[2634];
				12'd2635	: data1 <= weights[2635];
				12'd2636	: data1 <= weights[2636];
				12'd2637	: data1 <= weights[2637];
				12'd2638	: data1 <= weights[2638];
				12'd2639	: data1 <= weights[2639];
				12'd2640	: data1 <= weights[2640];
				12'd2641	: data1 <= weights[2641];
				12'd2642	: data1 <= weights[2642];
				12'd2643	: data1 <= weights[2643];
				12'd2644	: data1 <= weights[2644];
				12'd2645	: data1 <= weights[2645];
				12'd2646	: data1 <= weights[2646];
				12'd2647	: data1 <= weights[2647];
				12'd2648	: data1 <= weights[2648];
				12'd2649	: data1 <= weights[2649];
				12'd2650	: data1 <= weights[2650];
				12'd2651	: data1 <= weights[2651];
				12'd2652	: data1 <= weights[2652];
				12'd2653	: data1 <= weights[2653];
				12'd2654	: data1 <= weights[2654];
				12'd2655	: data1 <= weights[2655];
				12'd2656	: data1 <= weights[2656];
				12'd2657	: data1 <= weights[2657];
				12'd2658	: data1 <= weights[2658];
				12'd2659	: data1 <= weights[2659];
				12'd2660	: data1 <= weights[2660];
				12'd2661	: data1 <= weights[2661];
				12'd2662	: data1 <= weights[2662];
				12'd2663	: data1 <= weights[2663];
				12'd2664	: data1 <= weights[2664];
				12'd2665	: data1 <= weights[2665];
				12'd2666	: data1 <= weights[2666];
				12'd2667	: data1 <= weights[2667];
				12'd2668	: data1 <= weights[2668];
				12'd2669	: data1 <= weights[2669];
				12'd2670	: data1 <= weights[2670];
				12'd2671	: data1 <= weights[2671];
				12'd2672	: data1 <= weights[2672];
				12'd2673	: data1 <= weights[2673];
				12'd2674	: data1 <= weights[2674];
				12'd2675	: data1 <= weights[2675];
				12'd2676	: data1 <= weights[2676];
				12'd2677	: data1 <= weights[2677];
				12'd2678	: data1 <= weights[2678];
				12'd2679	: data1 <= weights[2679];
				12'd2680	: data1 <= weights[2680];
				12'd2681	: data1 <= weights[2681];
				12'd2682	: data1 <= weights[2682];
				12'd2683	: data1 <= weights[2683];
				12'd2684	: data1 <= weights[2684];
				12'd2685	: data1 <= weights[2685];
				12'd2686	: data1 <= weights[2686];
				12'd2687	: data1 <= weights[2687];
				12'd2688	: data1 <= weights[2688];
				12'd2689	: data1 <= weights[2689];
				12'd2690	: data1 <= weights[2690];
				12'd2691	: data1 <= weights[2691];
				12'd2692	: data1 <= weights[2692];
				12'd2693	: data1 <= weights[2693];
				12'd2694	: data1 <= weights[2694];
				12'd2695	: data1 <= weights[2695];
				12'd2696	: data1 <= weights[2696];
				12'd2697	: data1 <= weights[2697];
				12'd2698	: data1 <= weights[2698];
				12'd2699	: data1 <= weights[2699];
				12'd2700	: data1 <= weights[2700];
				12'd2701	: data1 <= weights[2701];
				12'd2702	: data1 <= weights[2702];
				12'd2703	: data1 <= weights[2703];
				12'd2704	: data1 <= weights[2704];
				12'd2705	: data1 <= weights[2705];
				12'd2706	: data1 <= weights[2706];
				12'd2707	: data1 <= weights[2707];
				12'd2708	: data1 <= weights[2708];
				12'd2709	: data1 <= weights[2709];
				12'd2710	: data1 <= weights[2710];
				12'd2711	: data1 <= weights[2711];
				12'd2712	: data1 <= weights[2712];
				12'd2713	: data1 <= weights[2713];
				12'd2714	: data1 <= weights[2714];
				12'd2715	: data1 <= weights[2715];
				12'd2716	: data1 <= weights[2716];
				12'd2717	: data1 <= weights[2717];
				12'd2718	: data1 <= weights[2718];
				12'd2719	: data1 <= weights[2719];
				12'd2720	: data1 <= weights[2720];
				12'd2721	: data1 <= weights[2721];
				12'd2722	: data1 <= weights[2722];
				12'd2723	: data1 <= weights[2723];
				12'd2724	: data1 <= weights[2724];
				12'd2725	: data1 <= weights[2725];
				12'd2726	: data1 <= weights[2726];
				12'd2727	: data1 <= weights[2727];
				12'd2728	: data1 <= weights[2728];
				12'd2729	: data1 <= weights[2729];
				12'd2730	: data1 <= weights[2730];
				12'd2731	: data1 <= weights[2731];
				12'd2732	: data1 <= weights[2732];
				12'd2733	: data1 <= weights[2733];
				12'd2734	: data1 <= weights[2734];
				12'd2735	: data1 <= weights[2735];
				12'd2736	: data1 <= weights[2736];
				12'd2737	: data1 <= weights[2737];
				12'd2738	: data1 <= weights[2738];
				12'd2739	: data1 <= weights[2739];
				12'd2740	: data1 <= weights[2740];
				12'd2741	: data1 <= weights[2741];
				12'd2742	: data1 <= weights[2742];
				12'd2743	: data1 <= weights[2743];
				12'd2744	: data1 <= weights[2744];
				12'd2745	: data1 <= weights[2745];
				12'd2746	: data1 <= weights[2746];
				12'd2747	: data1 <= weights[2747];
				12'd2748	: data1 <= weights[2748];
				12'd2749	: data1 <= weights[2749];
				12'd2750	: data1 <= weights[2750];
				12'd2751	: data1 <= weights[2751];
				12'd2752	: data1 <= weights[2752];
				12'd2753	: data1 <= weights[2753];
				12'd2754	: data1 <= weights[2754];
				12'd2755	: data1 <= weights[2755];
				12'd2756	: data1 <= weights[2756];
				12'd2757	: data1 <= weights[2757];
				12'd2758	: data1 <= weights[2758];
				12'd2759	: data1 <= weights[2759];
				12'd2760	: data1 <= weights[2760];
				12'd2761	: data1 <= weights[2761];
				12'd2762	: data1 <= weights[2762];
				12'd2763	: data1 <= weights[2763];
				12'd2764	: data1 <= weights[2764];
				12'd2765	: data1 <= weights[2765];
				12'd2766	: data1 <= weights[2766];
				12'd2767	: data1 <= weights[2767];
				12'd2768	: data1 <= weights[2768];
				12'd2769	: data1 <= weights[2769];
				12'd2770	: data1 <= weights[2770];
				12'd2771	: data1 <= weights[2771];
				12'd2772	: data1 <= weights[2772];
				12'd2773	: data1 <= weights[2773];
				12'd2774	: data1 <= weights[2774];
				12'd2775	: data1 <= weights[2775];
				12'd2776	: data1 <= weights[2776];
				12'd2777	: data1 <= weights[2777];
				12'd2778	: data1 <= weights[2778];
				12'd2779	: data1 <= weights[2779];
				12'd2780	: data1 <= weights[2780];
				12'd2781	: data1 <= weights[2781];
				12'd2782	: data1 <= weights[2782];
				12'd2783	: data1 <= weights[2783];
				12'd2784	: data1 <= weights[2784];
				12'd2785	: data1 <= weights[2785];
				12'd2786	: data1 <= weights[2786];
				12'd2787	: data1 <= weights[2787];
				12'd2788	: data1 <= weights[2788];
				12'd2789	: data1 <= weights[2789];
				12'd2790	: data1 <= weights[2790];
				12'd2791	: data1 <= weights[2791];
				12'd2792	: data1 <= weights[2792];
				12'd2793	: data1 <= weights[2793];
				12'd2794	: data1 <= weights[2794];
				12'd2795	: data1 <= weights[2795];
				12'd2796	: data1 <= weights[2796];
				12'd2797	: data1 <= weights[2797];
				12'd2798	: data1 <= weights[2798];
				12'd2799	: data1 <= weights[2799];
				12'd2800	: data1 <= weights[2800];
				12'd2801	: data1 <= weights[2801];
				12'd2802	: data1 <= weights[2802];
				12'd2803	: data1 <= weights[2803];
				12'd2804	: data1 <= weights[2804];
				12'd2805	: data1 <= weights[2805];
				12'd2806	: data1 <= weights[2806];
				12'd2807	: data1 <= weights[2807];
				12'd2808	: data1 <= weights[2808];
				12'd2809	: data1 <= weights[2809];
				12'd2810	: data1 <= weights[2810];
				12'd2811	: data1 <= weights[2811];
				12'd2812	: data1 <= weights[2812];
				12'd2813	: data1 <= weights[2813];
				12'd2814	: data1 <= weights[2814];
				12'd2815	: data1 <= weights[2815];
				12'd2816	: data1 <= weights[2816];
				12'd2817	: data1 <= weights[2817];
				12'd2818	: data1 <= weights[2818];
				12'd2819	: data1 <= weights[2819];
				12'd2820	: data1 <= weights[2820];
				12'd2821	: data1 <= weights[2821];
				12'd2822	: data1 <= weights[2822];
				12'd2823	: data1 <= weights[2823];
				12'd2824	: data1 <= weights[2824];
				12'd2825	: data1 <= weights[2825];
				12'd2826	: data1 <= weights[2826];
				12'd2827	: data1 <= weights[2827];
				12'd2828	: data1 <= weights[2828];
				12'd2829	: data1 <= weights[2829];
				12'd2830	: data1 <= weights[2830];
				12'd2831	: data1 <= weights[2831];
				12'd2832	: data1 <= weights[2832];
				12'd2833	: data1 <= weights[2833];
				12'd2834	: data1 <= weights[2834];
				12'd2835	: data1 <= weights[2835];
				12'd2836	: data1 <= weights[2836];
				12'd2837	: data1 <= weights[2837];
				12'd2838	: data1 <= weights[2838];
				12'd2839	: data1 <= weights[2839];
				12'd2840	: data1 <= weights[2840];
				12'd2841	: data1 <= weights[2841];
				12'd2842	: data1 <= weights[2842];
				12'd2843	: data1 <= weights[2843];
				12'd2844	: data1 <= weights[2844];
				12'd2845	: data1 <= weights[2845];
				12'd2846	: data1 <= weights[2846];
				12'd2847	: data1 <= weights[2847];
				12'd2848	: data1 <= weights[2848];
				12'd2849	: data1 <= weights[2849];
				12'd2850	: data1 <= weights[2850];
				12'd2851	: data1 <= weights[2851];
				12'd2852	: data1 <= weights[2852];
				12'd2853	: data1 <= weights[2853];
				12'd2854	: data1 <= weights[2854];
				12'd2855	: data1 <= weights[2855];
				12'd2856	: data1 <= weights[2856];
				12'd2857	: data1 <= weights[2857];
				12'd2858	: data1 <= weights[2858];
				12'd2859	: data1 <= weights[2859];
				12'd2860	: data1 <= weights[2860];
				12'd2861	: data1 <= weights[2861];
				12'd2862	: data1 <= weights[2862];
				12'd2863	: data1 <= weights[2863];
				12'd2864	: data1 <= weights[2864];
				12'd2865	: data1 <= weights[2865];
				12'd2866	: data1 <= weights[2866];
				12'd2867	: data1 <= weights[2867];
				12'd2868	: data1 <= weights[2868];
				12'd2869	: data1 <= weights[2869];
				12'd2870	: data1 <= weights[2870];
				12'd2871	: data1 <= weights[2871];
				12'd2872	: data1 <= weights[2872];
				12'd2873	: data1 <= weights[2873];
				12'd2874	: data1 <= weights[2874];
				12'd2875	: data1 <= weights[2875];
				12'd2876	: data1 <= weights[2876];
				12'd2877	: data1 <= weights[2877];
				12'd2878	: data1 <= weights[2878];
				12'd2879	: data1 <= weights[2879];
				12'd2880	: data1 <= weights[2880];
				12'd2881	: data1 <= weights[2881];
				12'd2882	: data1 <= weights[2882];
				12'd2883	: data1 <= weights[2883];
				12'd2884	: data1 <= weights[2884];
				12'd2885	: data1 <= weights[2885];
				12'd2886	: data1 <= weights[2886];
				12'd2887	: data1 <= weights[2887];
				12'd2888	: data1 <= weights[2888];
				12'd2889	: data1 <= weights[2889];
				12'd2890	: data1 <= weights[2890];
				12'd2891	: data1 <= weights[2891];
				12'd2892	: data1 <= weights[2892];
				12'd2893	: data1 <= weights[2893];
				12'd2894	: data1 <= weights[2894];
				12'd2895	: data1 <= weights[2895];
				12'd2896	: data1 <= weights[2896];
				12'd2897	: data1 <= weights[2897];
				12'd2898	: data1 <= weights[2898];
				12'd2899	: data1 <= weights[2899];
				12'd2900	: data1 <= weights[2900];
				12'd2901	: data1 <= weights[2901];
				12'd2902	: data1 <= weights[2902];
				12'd2903	: data1 <= weights[2903];
				12'd2904	: data1 <= weights[2904];
				12'd2905	: data1 <= weights[2905];
				12'd2906	: data1 <= weights[2906];
				12'd2907	: data1 <= weights[2907];
				12'd2908	: data1 <= weights[2908];
				12'd2909	: data1 <= weights[2909];
				12'd2910	: data1 <= weights[2910];
				12'd2911	: data1 <= weights[2911];
				12'd2912	: data1 <= weights[2912];
				12'd2913	: data1 <= weights[2913];
				12'd2914	: data1 <= weights[2914];
				12'd2915	: data1 <= weights[2915];
				12'd2916	: data1 <= weights[2916];
				12'd2917	: data1 <= weights[2917];
				12'd2918	: data1 <= weights[2918];
				12'd2919	: data1 <= weights[2919];
				12'd2920	: data1 <= weights[2920];
				12'd2921	: data1 <= weights[2921];
				12'd2922	: data1 <= weights[2922];
				12'd2923	: data1 <= weights[2923];
				12'd2924	: data1 <= weights[2924];
				12'd2925	: data1 <= weights[2925];
				12'd2926	: data1 <= weights[2926];
				12'd2927	: data1 <= weights[2927];
				12'd2928	: data1 <= weights[2928];
				12'd2929	: data1 <= weights[2929];
				12'd2930	: data1 <= weights[2930];
				12'd2931	: data1 <= weights[2931];
				12'd2932	: data1 <= weights[2932];
				12'd2933	: data1 <= weights[2933];
				12'd2934	: data1 <= weights[2934];
				12'd2935	: data1 <= weights[2935];
				12'd2936	: data1 <= weights[2936];
				12'd2937	: data1 <= weights[2937];
				12'd2938	: data1 <= weights[2938];
				12'd2939	: data1 <= weights[2939];
				12'd2940	: data1 <= weights[2940];
				12'd2941	: data1 <= weights[2941];
				12'd2942	: data1 <= weights[2942];
				12'd2943	: data1 <= weights[2943];
				12'd2944	: data1 <= weights[2944];
				12'd2945	: data1 <= weights[2945];
				12'd2946	: data1 <= weights[2946];
				12'd2947	: data1 <= weights[2947];
				12'd2948	: data1 <= weights[2948];
				12'd2949	: data1 <= weights[2949];
				12'd2950	: data1 <= weights[2950];
				12'd2951	: data1 <= weights[2951];
				12'd2952	: data1 <= weights[2952];
				12'd2953	: data1 <= weights[2953];
				12'd2954	: data1 <= weights[2954];
				12'd2955	: data1 <= weights[2955];
				12'd2956	: data1 <= weights[2956];
				12'd2957	: data1 <= weights[2957];
				12'd2958	: data1 <= weights[2958];
				12'd2959	: data1 <= weights[2959];
				12'd2960	: data1 <= weights[2960];
				12'd2961	: data1 <= weights[2961];
				12'd2962	: data1 <= weights[2962];
				12'd2963	: data1 <= weights[2963];
				12'd2964	: data1 <= weights[2964];
				12'd2965	: data1 <= weights[2965];
				12'd2966	: data1 <= weights[2966];
				12'd2967	: data1 <= weights[2967];
				12'd2968	: data1 <= weights[2968];
				12'd2969	: data1 <= weights[2969];
				12'd2970	: data1 <= weights[2970];
				12'd2971	: data1 <= weights[2971];
				12'd2972	: data1 <= weights[2972];
				12'd2973	: data1 <= weights[2973];
				12'd2974	: data1 <= weights[2974];
				12'd2975	: data1 <= weights[2975];
				12'd2976	: data1 <= weights[2976];
				12'd2977	: data1 <= weights[2977];
				12'd2978	: data1 <= weights[2978];
				12'd2979	: data1 <= weights[2979];
				12'd2980	: data1 <= weights[2980];
				12'd2981	: data1 <= weights[2981];
				12'd2982	: data1 <= weights[2982];
				12'd2983	: data1 <= weights[2983];
				12'd2984	: data1 <= weights[2984];
				12'd2985	: data1 <= weights[2985];
				12'd2986	: data1 <= weights[2986];
				12'd2987	: data1 <= weights[2987];
				12'd2988	: data1 <= weights[2988];
				12'd2989	: data1 <= weights[2989];
				12'd2990	: data1 <= weights[2990];
				12'd2991	: data1 <= weights[2991];
				12'd2992	: data1 <= weights[2992];
				12'd2993	: data1 <= weights[2993];
				12'd2994	: data1 <= weights[2994];
				12'd2995	: data1 <= weights[2995];
				12'd2996	: data1 <= weights[2996];
				12'd2997	: data1 <= weights[2997];
				12'd2998	: data1 <= weights[2998];
				12'd2999	: data1 <= weights[2999];
				12'd3000	: data1 <= weights[3000];
				12'd3001	: data1 <= weights[3001];
				12'd3002	: data1 <= weights[3002];
				12'd3003	: data1 <= weights[3003];
				12'd3004	: data1 <= weights[3004];
				12'd3005	: data1 <= weights[3005];
				12'd3006	: data1 <= weights[3006];
				12'd3007	: data1 <= weights[3007];
				12'd3008	: data1 <= weights[3008];
				12'd3009	: data1 <= weights[3009];
				12'd3010	: data1 <= weights[3010];
				12'd3011	: data1 <= weights[3011];
				12'd3012	: data1 <= weights[3012];
				12'd3013	: data1 <= weights[3013];
				12'd3014	: data1 <= weights[3014];
				12'd3015	: data1 <= weights[3015];
				12'd3016	: data1 <= weights[3016];
				12'd3017	: data1 <= weights[3017];
				12'd3018	: data1 <= weights[3018];
				12'd3019	: data1 <= weights[3019];
				12'd3020	: data1 <= weights[3020];
				12'd3021	: data1 <= weights[3021];
				12'd3022	: data1 <= weights[3022];
				12'd3023	: data1 <= weights[3023];
				12'd3024	: data1 <= weights[3024];
				12'd3025	: data1 <= weights[3025];
				12'd3026	: data1 <= weights[3026];
				12'd3027	: data1 <= weights[3027];
				12'd3028	: data1 <= weights[3028];
				12'd3029	: data1 <= weights[3029];
				12'd3030	: data1 <= weights[3030];
				12'd3031	: data1 <= weights[3031];
				12'd3032	: data1 <= weights[3032];
				12'd3033	: data1 <= weights[3033];
				12'd3034	: data1 <= weights[3034];
				12'd3035	: data1 <= weights[3035];
				12'd3036	: data1 <= weights[3036];
				12'd3037	: data1 <= weights[3037];
				12'd3038	: data1 <= weights[3038];
				12'd3039	: data1 <= weights[3039];
				12'd3040	: data1 <= weights[3040];
				12'd3041	: data1 <= weights[3041];
				12'd3042	: data1 <= weights[3042];
				12'd3043	: data1 <= weights[3043];
				12'd3044	: data1 <= weights[3044];
				12'd3045	: data1 <= weights[3045];
				12'd3046	: data1 <= weights[3046];
				12'd3047	: data1 <= weights[3047];
				12'd3048	: data1 <= weights[3048];
				12'd3049	: data1 <= weights[3049];
				12'd3050	: data1 <= weights[3050];
				12'd3051	: data1 <= weights[3051];
				12'd3052	: data1 <= weights[3052];
				12'd3053	: data1 <= weights[3053];
				12'd3054	: data1 <= weights[3054];
				12'd3055	: data1 <= weights[3055];
				12'd3056	: data1 <= weights[3056];
				12'd3057	: data1 <= weights[3057];
				12'd3058	: data1 <= weights[3058];
				12'd3059	: data1 <= weights[3059];
				12'd3060	: data1 <= weights[3060];
				12'd3061	: data1 <= weights[3061];
				12'd3062	: data1 <= weights[3062];
				12'd3063	: data1 <= weights[3063];
				12'd3064	: data1 <= weights[3064];
				12'd3065	: data1 <= weights[3065];
				12'd3066	: data1 <= weights[3066];
				12'd3067	: data1 <= weights[3067];
				12'd3068	: data1 <= weights[3068];
				12'd3069	: data1 <= weights[3069];
				12'd3070	: data1 <= weights[3070];
				12'd3071	: data1 <= weights[3071];
				12'd3072	: data1 <= weights[3072];
				12'd3073	: data1 <= weights[3073];
				12'd3074	: data1 <= weights[3074];
				12'd3075	: data1 <= weights[3075];
				12'd3076	: data1 <= weights[3076];
				12'd3077	: data1 <= weights[3077];
				12'd3078	: data1 <= weights[3078];
				12'd3079	: data1 <= weights[3079];
				12'd3080	: data1 <= weights[3080];
				12'd3081	: data1 <= weights[3081];
				12'd3082	: data1 <= weights[3082];
				12'd3083	: data1 <= weights[3083];
				12'd3084	: data1 <= weights[3084];
				12'd3085	: data1 <= weights[3085];
				12'd3086	: data1 <= weights[3086];
				12'd3087	: data1 <= weights[3087];
				12'd3088	: data1 <= weights[3088];
				12'd3089	: data1 <= weights[3089];
				12'd3090	: data1 <= weights[3090];
				12'd3091	: data1 <= weights[3091];
				12'd3092	: data1 <= weights[3092];
				12'd3093	: data1 <= weights[3093];
				12'd3094	: data1 <= weights[3094];
				12'd3095	: data1 <= weights[3095];
				12'd3096	: data1 <= weights[3096];
				12'd3097	: data1 <= weights[3097];
				12'd3098	: data1 <= weights[3098];
				12'd3099	: data1 <= weights[3099];
				12'd3100	: data1 <= weights[3100];
				12'd3101	: data1 <= weights[3101];
				12'd3102	: data1 <= weights[3102];
				12'd3103	: data1 <= weights[3103];
				12'd3104	: data1 <= weights[3104];
				12'd3105	: data1 <= weights[3105];
				12'd3106	: data1 <= weights[3106];
				12'd3107	: data1 <= weights[3107];
				12'd3108	: data1 <= weights[3108];
				12'd3109	: data1 <= weights[3109];
				12'd3110	: data1 <= weights[3110];
				12'd3111	: data1 <= weights[3111];
				12'd3112	: data1 <= weights[3112];
				12'd3113	: data1 <= weights[3113];
				12'd3114	: data1 <= weights[3114];
				12'd3115	: data1 <= weights[3115];
				12'd3116	: data1 <= weights[3116];
				12'd3117	: data1 <= weights[3117];
				12'd3118	: data1 <= weights[3118];
				12'd3119	: data1 <= weights[3119];
				12'd3120	: data1 <= weights[3120];
				12'd3121	: data1 <= weights[3121];
				12'd3122	: data1 <= weights[3122];
				12'd3123	: data1 <= weights[3123];
				12'd3124	: data1 <= weights[3124];
				12'd3125	: data1 <= weights[3125];
				12'd3126	: data1 <= weights[3126];
				12'd3127	: data1 <= weights[3127];
				12'd3128	: data1 <= weights[3128];
				12'd3129	: data1 <= weights[3129];
				12'd3130	: data1 <= weights[3130];
				12'd3131	: data1 <= weights[3131];
				12'd3132	: data1 <= weights[3132];
				12'd3133	: data1 <= weights[3133];
				12'd3134	: data1 <= weights[3134];
				12'd3135	: data1 <= weights[3135];
				12'd3136	: data1 <= weights[3136];
				12'd3137	: data1 <= weights[3137];
				12'd3138	: data1 <= weights[3138];
				12'd3139	: data1 <= weights[3139];
				12'd3140	: data1 <= weights[3140];
				12'd3141	: data1 <= weights[3141];
				12'd3142	: data1 <= weights[3142];
				12'd3143	: data1 <= weights[3143];
				12'd3144	: data1 <= weights[3144];
				12'd3145	: data1 <= weights[3145];
				12'd3146	: data1 <= weights[3146];
				12'd3147	: data1 <= weights[3147];
				12'd3148	: data1 <= weights[3148];
				12'd3149	: data1 <= weights[3149];
				12'd3150	: data1 <= weights[3150];
				12'd3151	: data1 <= weights[3151];
				12'd3152	: data1 <= weights[3152];
				12'd3153	: data1 <= weights[3153];
				12'd3154	: data1 <= weights[3154];
				12'd3155	: data1 <= weights[3155];
				12'd3156	: data1 <= weights[3156];
				12'd3157	: data1 <= weights[3157];
				12'd3158	: data1 <= weights[3158];
				12'd3159	: data1 <= weights[3159];
				12'd3160	: data1 <= weights[3160];
				12'd3161	: data1 <= weights[3161];
				12'd3162	: data1 <= weights[3162];
				12'd3163	: data1 <= weights[3163];
				12'd3164	: data1 <= weights[3164];
				12'd3165	: data1 <= weights[3165];
				12'd3166	: data1 <= weights[3166];
				12'd3167	: data1 <= weights[3167];
				12'd3168	: data1 <= weights[3168];
				12'd3169	: data1 <= weights[3169];
				12'd3170	: data1 <= weights[3170];
				12'd3171	: data1 <= weights[3171];
				12'd3172	: data1 <= weights[3172];
				12'd3173	: data1 <= weights[3173];
				12'd3174	: data1 <= weights[3174];
				12'd3175	: data1 <= weights[3175];
				12'd3176	: data1 <= weights[3176];
				12'd3177	: data1 <= weights[3177];
				12'd3178	: data1 <= weights[3178];
				12'd3179	: data1 <= weights[3179];
				12'd3180	: data1 <= weights[3180];
				12'd3181	: data1 <= weights[3181];
				12'd3182	: data1 <= weights[3182];
				12'd3183	: data1 <= weights[3183];
				12'd3184	: data1 <= weights[3184];
				12'd3185	: data1 <= weights[3185];
				12'd3186	: data1 <= weights[3186];
				12'd3187	: data1 <= weights[3187];
				12'd3188	: data1 <= weights[3188];
				12'd3189	: data1 <= weights[3189];
				12'd3190	: data1 <= weights[3190];
				12'd3191	: data1 <= weights[3191];
				12'd3192	: data1 <= weights[3192];
				12'd3193	: data1 <= weights[3193];
				12'd3194	: data1 <= weights[3194];
				12'd3195	: data1 <= weights[3195];
				12'd3196	: data1 <= weights[3196];
				12'd3197	: data1 <= weights[3197];
				12'd3198	: data1 <= weights[3198];
				12'd3199	: data1 <= weights[3199];
				12'd3200	: data1 <= weights[3200];
				12'd3201	: data1 <= weights[3201];
				12'd3202	: data1 <= weights[3202];
				12'd3203	: data1 <= weights[3203];
				12'd3204	: data1 <= weights[3204];
				12'd3205	: data1 <= weights[3205];
				12'd3206	: data1 <= weights[3206];
				12'd3207	: data1 <= weights[3207];
				12'd3208	: data1 <= weights[3208];
				12'd3209	: data1 <= weights[3209];
				12'd3210	: data1 <= weights[3210];
				12'd3211	: data1 <= weights[3211];
				12'd3212	: data1 <= weights[3212];
				12'd3213	: data1 <= weights[3213];
				12'd3214	: data1 <= weights[3214];
				12'd3215	: data1 <= weights[3215];
				12'd3216	: data1 <= weights[3216];
				12'd3217	: data1 <= weights[3217];
				12'd3218	: data1 <= weights[3218];
				12'd3219	: data1 <= weights[3219];
				12'd3220	: data1 <= weights[3220];
				12'd3221	: data1 <= weights[3221];
				12'd3222	: data1 <= weights[3222];
				12'd3223	: data1 <= weights[3223];
				12'd3224	: data1 <= weights[3224];
				12'd3225	: data1 <= weights[3225];
				12'd3226	: data1 <= weights[3226];
				12'd3227	: data1 <= weights[3227];
				12'd3228	: data1 <= weights[3228];
				12'd3229	: data1 <= weights[3229];
				12'd3230	: data1 <= weights[3230];
				12'd3231	: data1 <= weights[3231];
				12'd3232	: data1 <= weights[3232];
				12'd3233	: data1 <= weights[3233];
				12'd3234	: data1 <= weights[3234];
				12'd3235	: data1 <= weights[3235];
				12'd3236	: data1 <= weights[3236];
				12'd3237	: data1 <= weights[3237];
				12'd3238	: data1 <= weights[3238];
				12'd3239	: data1 <= weights[3239];
				12'd3240	: data1 <= weights[3240];
				12'd3241	: data1 <= weights[3241];
				12'd3242	: data1 <= weights[3242];
				12'd3243	: data1 <= weights[3243];
				12'd3244	: data1 <= weights[3244];
				12'd3245	: data1 <= weights[3245];
				12'd3246	: data1 <= weights[3246];
				12'd3247	: data1 <= weights[3247];
				12'd3248	: data1 <= weights[3248];
				12'd3249	: data1 <= weights[3249];
				12'd3250	: data1 <= weights[3250];
				12'd3251	: data1 <= weights[3251];
				12'd3252	: data1 <= weights[3252];
				12'd3253	: data1 <= weights[3253];
				12'd3254	: data1 <= weights[3254];
				12'd3255	: data1 <= weights[3255];
				12'd3256	: data1 <= weights[3256];
				12'd3257	: data1 <= weights[3257];
				12'd3258	: data1 <= weights[3258];
				12'd3259	: data1 <= weights[3259];
				12'd3260	: data1 <= weights[3260];
				12'd3261	: data1 <= weights[3261];
				12'd3262	: data1 <= weights[3262];
				12'd3263	: data1 <= weights[3263];
				12'd3264	: data1 <= weights[3264];
				12'd3265	: data1 <= weights[3265];
				12'd3266	: data1 <= weights[3266];
				12'd3267	: data1 <= weights[3267];
				12'd3268	: data1 <= weights[3268];
				12'd3269	: data1 <= weights[3269];
				12'd3270	: data1 <= weights[3270];
				12'd3271	: data1 <= weights[3271];
				12'd3272	: data1 <= weights[3272];
				12'd3273	: data1 <= weights[3273];
				12'd3274	: data1 <= weights[3274];
				12'd3275	: data1 <= weights[3275];
				12'd3276	: data1 <= weights[3276];
				12'd3277	: data1 <= weights[3277];
				12'd3278	: data1 <= weights[3278];
				12'd3279	: data1 <= weights[3279];
				12'd3280	: data1 <= weights[3280];
				12'd3281	: data1 <= weights[3281];
				12'd3282	: data1 <= weights[3282];
				12'd3283	: data1 <= weights[3283];
				12'd3284	: data1 <= weights[3284];
				12'd3285	: data1 <= weights[3285];
				12'd3286	: data1 <= weights[3286];
				12'd3287	: data1 <= weights[3287];
				12'd3288	: data1 <= weights[3288];
				12'd3289	: data1 <= weights[3289];
				12'd3290	: data1 <= weights[3290];
				12'd3291	: data1 <= weights[3291];
				12'd3292	: data1 <= weights[3292];
				12'd3293	: data1 <= weights[3293];
				12'd3294	: data1 <= weights[3294];
				12'd3295	: data1 <= weights[3295];
				12'd3296	: data1 <= weights[3296];
				12'd3297	: data1 <= weights[3297];
				12'd3298	: data1 <= weights[3298];
				12'd3299	: data1 <= weights[3299];
				12'd3300	: data1 <= weights[3300];
				12'd3301	: data1 <= weights[3301];
				12'd3302	: data1 <= weights[3302];
				12'd3303	: data1 <= weights[3303];
				12'd3304	: data1 <= weights[3304];
				12'd3305	: data1 <= weights[3305];
				12'd3306	: data1 <= weights[3306];
				12'd3307	: data1 <= weights[3307];
				12'd3308	: data1 <= weights[3308];
				12'd3309	: data1 <= weights[3309];
				12'd3310	: data1 <= weights[3310];
				12'd3311	: data1 <= weights[3311];
				12'd3312	: data1 <= weights[3312];
				12'd3313	: data1 <= weights[3313];
				12'd3314	: data1 <= weights[3314];
				12'd3315	: data1 <= weights[3315];
				12'd3316	: data1 <= weights[3316];
				12'd3317	: data1 <= weights[3317];
				12'd3318	: data1 <= weights[3318];
				12'd3319	: data1 <= weights[3319];
				12'd3320	: data1 <= weights[3320];
				12'd3321	: data1 <= weights[3321];
				12'd3322	: data1 <= weights[3322];
				12'd3323	: data1 <= weights[3323];
				12'd3324	: data1 <= weights[3324];
				12'd3325	: data1 <= weights[3325];
				12'd3326	: data1 <= weights[3326];
				12'd3327	: data1 <= weights[3327];
				12'd3328	: data1 <= weights[3328];
				12'd3329	: data1 <= weights[3329];
				12'd3330	: data1 <= weights[3330];
				12'd3331	: data1 <= weights[3331];
				12'd3332	: data1 <= weights[3332];
				12'd3333	: data1 <= weights[3333];
				12'd3334	: data1 <= weights[3334];
				12'd3335	: data1 <= weights[3335];
				12'd3336	: data1 <= weights[3336];
				12'd3337	: data1 <= weights[3337];
				12'd3338	: data1 <= weights[3338];
				12'd3339	: data1 <= weights[3339];
				12'd3340	: data1 <= weights[3340];
				12'd3341	: data1 <= weights[3341];
				12'd3342	: data1 <= weights[3342];
				12'd3343	: data1 <= weights[3343];
				12'd3344	: data1 <= weights[3344];
				12'd3345	: data1 <= weights[3345];
				12'd3346	: data1 <= weights[3346];
				12'd3347	: data1 <= weights[3347];
				12'd3348	: data1 <= weights[3348];
				12'd3349	: data1 <= weights[3349];
				12'd3350	: data1 <= weights[3350];
				12'd3351	: data1 <= weights[3351];
				12'd3352	: data1 <= weights[3352];
				12'd3353	: data1 <= weights[3353];
				12'd3354	: data1 <= weights[3354];
				12'd3355	: data1 <= weights[3355];
				12'd3356	: data1 <= weights[3356];
				12'd3357	: data1 <= weights[3357];
				12'd3358	: data1 <= weights[3358];
				12'd3359	: data1 <= weights[3359];
				12'd3360	: data1 <= weights[3360];
				12'd3361	: data1 <= weights[3361];
				12'd3362	: data1 <= weights[3362];
				12'd3363	: data1 <= weights[3363];
				12'd3364	: data1 <= weights[3364];
				12'd3365	: data1 <= weights[3365];
				12'd3366	: data1 <= weights[3366];
				12'd3367	: data1 <= weights[3367];
				12'd3368	: data1 <= weights[3368];
				12'd3369	: data1 <= weights[3369];
				12'd3370	: data1 <= weights[3370];
				12'd3371	: data1 <= weights[3371];
				12'd3372	: data1 <= weights[3372];
				12'd3373	: data1 <= weights[3373];
				12'd3374	: data1 <= weights[3374];
				12'd3375	: data1 <= weights[3375];
				12'd3376	: data1 <= weights[3376];
				12'd3377	: data1 <= weights[3377];
				12'd3378	: data1 <= weights[3378];
				12'd3379	: data1 <= weights[3379];
				12'd3380	: data1 <= weights[3380];
				12'd3381	: data1 <= weights[3381];
				12'd3382	: data1 <= weights[3382];
				12'd3383	: data1 <= weights[3383];
				12'd3384	: data1 <= weights[3384];
				12'd3385	: data1 <= weights[3385];
				12'd3386	: data1 <= weights[3386];
				12'd3387	: data1 <= weights[3387];
				12'd3388	: data1 <= weights[3388];
				12'd3389	: data1 <= weights[3389];
				12'd3390	: data1 <= weights[3390];
				12'd3391	: data1 <= weights[3391];
				12'd3392	: data1 <= weights[3392];
				12'd3393	: data1 <= weights[3393];
				12'd3394	: data1 <= weights[3394];
				12'd3395	: data1 <= weights[3395];
				12'd3396	: data1 <= weights[3396];
				12'd3397	: data1 <= weights[3397];
				12'd3398	: data1 <= weights[3398];
				12'd3399	: data1 <= weights[3399];
				12'd3400	: data1 <= weights[3400];
				12'd3401	: data1 <= weights[3401];
				12'd3402	: data1 <= weights[3402];
				12'd3403	: data1 <= weights[3403];
				12'd3404	: data1 <= weights[3404];
				12'd3405	: data1 <= weights[3405];
				12'd3406	: data1 <= weights[3406];
				12'd3407	: data1 <= weights[3407];
				12'd3408	: data1 <= weights[3408];
				12'd3409	: data1 <= weights[3409];
				12'd3410	: data1 <= weights[3410];
				12'd3411	: data1 <= weights[3411];
				12'd3412	: data1 <= weights[3412];
				12'd3413	: data1 <= weights[3413];
				12'd3414	: data1 <= weights[3414];
				12'd3415	: data1 <= weights[3415];
				12'd3416	: data1 <= weights[3416];
				12'd3417	: data1 <= weights[3417];
				12'd3418	: data1 <= weights[3418];
				12'd3419	: data1 <= weights[3419];
				12'd3420	: data1 <= weights[3420];
				12'd3421	: data1 <= weights[3421];
				12'd3422	: data1 <= weights[3422];
				12'd3423	: data1 <= weights[3423];
				12'd3424	: data1 <= weights[3424];
				12'd3425	: data1 <= weights[3425];
				12'd3426	: data1 <= weights[3426];
				12'd3427	: data1 <= weights[3427];
				12'd3428	: data1 <= weights[3428];
				12'd3429	: data1 <= weights[3429];
				12'd3430	: data1 <= weights[3430];
				12'd3431	: data1 <= weights[3431];
				12'd3432	: data1 <= weights[3432];
				12'd3433	: data1 <= weights[3433];
				12'd3434	: data1 <= weights[3434];
				12'd3435	: data1 <= weights[3435];
				12'd3436	: data1 <= weights[3436];
				12'd3437	: data1 <= weights[3437];
				12'd3438	: data1 <= weights[3438];
				12'd3439	: data1 <= weights[3439];
				12'd3440	: data1 <= weights[3440];
				12'd3441	: data1 <= weights[3441];
				12'd3442	: data1 <= weights[3442];
				12'd3443	: data1 <= weights[3443];
				12'd3444	: data1 <= weights[3444];
				12'd3445	: data1 <= weights[3445];
				12'd3446	: data1 <= weights[3446];
				12'd3447	: data1 <= weights[3447];
				12'd3448	: data1 <= weights[3448];
				12'd3449	: data1 <= weights[3449];
				12'd3450	: data1 <= weights[3450];
				12'd3451	: data1 <= weights[3451];
				12'd3452	: data1 <= weights[3452];
				12'd3453	: data1 <= weights[3453];
				12'd3454	: data1 <= weights[3454];
				12'd3455	: data1 <= weights[3455];
				12'd3456	: data1 <= weights[3456];
				12'd3457	: data1 <= weights[3457];
				12'd3458	: data1 <= weights[3458];
				12'd3459	: data1 <= weights[3459];
				12'd3460	: data1 <= weights[3460];
				12'd3461	: data1 <= weights[3461];
				12'd3462	: data1 <= weights[3462];
				12'd3463	: data1 <= weights[3463];
				12'd3464	: data1 <= weights[3464];
				12'd3465	: data1 <= weights[3465];
				12'd3466	: data1 <= weights[3466];
				12'd3467	: data1 <= weights[3467];
				12'd3468	: data1 <= weights[3468];
				12'd3469	: data1 <= weights[3469];
				12'd3470	: data1 <= weights[3470];
				12'd3471	: data1 <= weights[3471];
				12'd3472	: data1 <= weights[3472];
				12'd3473	: data1 <= weights[3473];
				12'd3474	: data1 <= weights[3474];
				12'd3475	: data1 <= weights[3475];
				12'd3476	: data1 <= weights[3476];
				12'd3477	: data1 <= weights[3477];
				12'd3478	: data1 <= weights[3478];
				12'd3479	: data1 <= weights[3479];
				12'd3480	: data1 <= weights[3480];
				12'd3481	: data1 <= weights[3481];
				12'd3482	: data1 <= weights[3482];
				12'd3483	: data1 <= weights[3483];
				12'd3484	: data1 <= weights[3484];
				12'd3485	: data1 <= weights[3485];
				12'd3486	: data1 <= weights[3486];
				12'd3487	: data1 <= weights[3487];
				12'd3488	: data1 <= weights[3488];
				12'd3489	: data1 <= weights[3489];
				12'd3490	: data1 <= weights[3490];
				12'd3491	: data1 <= weights[3491];
				12'd3492	: data1 <= weights[3492];
				12'd3493	: data1 <= weights[3493];
				12'd3494	: data1 <= weights[3494];
				12'd3495	: data1 <= weights[3495];
				12'd3496	: data1 <= weights[3496];
				12'd3497	: data1 <= weights[3497];
				12'd3498	: data1 <= weights[3498];
				12'd3499	: data1 <= weights[3499];
				12'd3500	: data1 <= weights[3500];
				12'd3501	: data1 <= weights[3501];
				12'd3502	: data1 <= weights[3502];
				12'd3503	: data1 <= weights[3503];
				12'd3504	: data1 <= weights[3504];
				12'd3505	: data1 <= weights[3505];
				12'd3506	: data1 <= weights[3506];
				12'd3507	: data1 <= weights[3507];
				12'd3508	: data1 <= weights[3508];
				12'd3509	: data1 <= weights[3509];
				12'd3510	: data1 <= weights[3510];
				12'd3511	: data1 <= weights[3511];
				12'd3512	: data1 <= weights[3512];
				12'd3513	: data1 <= weights[3513];
				12'd3514	: data1 <= weights[3514];
				12'd3515	: data1 <= weights[3515];
				12'd3516	: data1 <= weights[3516];
				12'd3517	: data1 <= weights[3517];
				12'd3518	: data1 <= weights[3518];
				12'd3519	: data1 <= weights[3519];
				12'd3520	: data1 <= weights[3520];
				12'd3521	: data1 <= weights[3521];
				12'd3522	: data1 <= weights[3522];
				12'd3523	: data1 <= weights[3523];
				12'd3524	: data1 <= weights[3524];
				12'd3525	: data1 <= weights[3525];
				12'd3526	: data1 <= weights[3526];
				12'd3527	: data1 <= weights[3527];
				12'd3528	: data1 <= weights[3528];
				12'd3529	: data1 <= weights[3529];
				12'd3530	: data1 <= weights[3530];
				12'd3531	: data1 <= weights[3531];
				12'd3532	: data1 <= weights[3532];
				12'd3533	: data1 <= weights[3533];
				12'd3534	: data1 <= weights[3534];
				12'd3535	: data1 <= weights[3535];
				12'd3536	: data1 <= weights[3536];
				12'd3537	: data1 <= weights[3537];
				12'd3538	: data1 <= weights[3538];
				12'd3539	: data1 <= weights[3539];
				12'd3540	: data1 <= weights[3540];
				12'd3541	: data1 <= weights[3541];
				12'd3542	: data1 <= weights[3542];
				12'd3543	: data1 <= weights[3543];
				12'd3544	: data1 <= weights[3544];
				12'd3545	: data1 <= weights[3545];
				12'd3546	: data1 <= weights[3546];
				12'd3547	: data1 <= weights[3547];
				12'd3548	: data1 <= weights[3548];
				12'd3549	: data1 <= weights[3549];
				12'd3550	: data1 <= weights[3550];
				12'd3551	: data1 <= weights[3551];
				12'd3552	: data1 <= weights[3552];
				12'd3553	: data1 <= weights[3553];
				12'd3554	: data1 <= weights[3554];
				12'd3555	: data1 <= weights[3555];
				12'd3556	: data1 <= weights[3556];
				12'd3557	: data1 <= weights[3557];
				12'd3558	: data1 <= weights[3558];
				12'd3559	: data1 <= weights[3559];
				12'd3560	: data1 <= weights[3560];
				12'd3561	: data1 <= weights[3561];
				12'd3562	: data1 <= weights[3562];
				12'd3563	: data1 <= weights[3563];
				12'd3564	: data1 <= weights[3564];
				12'd3565	: data1 <= weights[3565];
				12'd3566	: data1 <= weights[3566];
				12'd3567	: data1 <= weights[3567];
				12'd3568	: data1 <= weights[3568];
				12'd3569	: data1 <= weights[3569];
				12'd3570	: data1 <= weights[3570];
				12'd3571	: data1 <= weights[3571];
				12'd3572	: data1 <= weights[3572];
				12'd3573	: data1 <= weights[3573];
				12'd3574	: data1 <= weights[3574];
				12'd3575	: data1 <= weights[3575];
				12'd3576	: data1 <= weights[3576];
				12'd3577	: data1 <= weights[3577];
				12'd3578	: data1 <= weights[3578];
				12'd3579	: data1 <= weights[3579];
				12'd3580	: data1 <= weights[3580];
				12'd3581	: data1 <= weights[3581];
				12'd3582	: data1 <= weights[3582];
				12'd3583	: data1 <= weights[3583];
				12'd3584	: data1 <= weights[3584];
				12'd3585	: data1 <= weights[3585];
				12'd3586	: data1 <= weights[3586];
				12'd3587	: data1 <= weights[3587];
				12'd3588	: data1 <= weights[3588];
				12'd3589	: data1 <= weights[3589];
				12'd3590	: data1 <= weights[3590];
				12'd3591	: data1 <= weights[3591];
				12'd3592	: data1 <= weights[3592];
				12'd3593	: data1 <= weights[3593];
				12'd3594	: data1 <= weights[3594];
				12'd3595	: data1 <= weights[3595];
				12'd3596	: data1 <= weights[3596];
				12'd3597	: data1 <= weights[3597];
				12'd3598	: data1 <= weights[3598];
				12'd3599	: data1 <= weights[3599];
				12'd3600	: data1 <= weights[3600];
				12'd3601	: data1 <= weights[3601];
				12'd3602	: data1 <= weights[3602];
				12'd3603	: data1 <= weights[3603];
				12'd3604	: data1 <= weights[3604];
				12'd3605	: data1 <= weights[3605];
				12'd3606	: data1 <= weights[3606];
				12'd3607	: data1 <= weights[3607];
				12'd3608	: data1 <= weights[3608];
				12'd3609	: data1 <= weights[3609];
				12'd3610	: data1 <= weights[3610];
				12'd3611	: data1 <= weights[3611];
				12'd3612	: data1 <= weights[3612];
				12'd3613	: data1 <= weights[3613];
				12'd3614	: data1 <= weights[3614];
				12'd3615	: data1 <= weights[3615];
				12'd3616	: data1 <= weights[3616];
				12'd3617	: data1 <= weights[3617];
				12'd3618	: data1 <= weights[3618];
				12'd3619	: data1 <= weights[3619];
				12'd3620	: data1 <= weights[3620];
				12'd3621	: data1 <= weights[3621];
				12'd3622	: data1 <= weights[3622];
				12'd3623	: data1 <= weights[3623];
				12'd3624	: data1 <= weights[3624];
				12'd3625	: data1 <= weights[3625];
				12'd3626	: data1 <= weights[3626];
				12'd3627	: data1 <= weights[3627];
				12'd3628	: data1 <= weights[3628];
				12'd3629	: data1 <= weights[3629];
				12'd3630	: data1 <= weights[3630];
				12'd3631	: data1 <= weights[3631];
				12'd3632	: data1 <= weights[3632];
				12'd3633	: data1 <= weights[3633];
				12'd3634	: data1 <= weights[3634];
				12'd3635	: data1 <= weights[3635];
				12'd3636	: data1 <= weights[3636];
				12'd3637	: data1 <= weights[3637];
				12'd3638	: data1 <= weights[3638];
				12'd3639	: data1 <= weights[3639];
				12'd3640	: data1 <= weights[3640];
				12'd3641	: data1 <= weights[3641];
				12'd3642	: data1 <= weights[3642];
				12'd3643	: data1 <= weights[3643];
				12'd3644	: data1 <= weights[3644];
				12'd3645	: data1 <= weights[3645];
				12'd3646	: data1 <= weights[3646];
				12'd3647	: data1 <= weights[3647];
				12'd3648	: data1 <= weights[3648];
				12'd3649	: data1 <= weights[3649];
				12'd3650	: data1 <= weights[3650];
				12'd3651	: data1 <= weights[3651];
				12'd3652	: data1 <= weights[3652];
				12'd3653	: data1 <= weights[3653];
				12'd3654	: data1 <= weights[3654];
				12'd3655	: data1 <= weights[3655];
				12'd3656	: data1 <= weights[3656];
				12'd3657	: data1 <= weights[3657];
				12'd3658	: data1 <= weights[3658];
				12'd3659	: data1 <= weights[3659];
				12'd3660	: data1 <= weights[3660];
				12'd3661	: data1 <= weights[3661];
				12'd3662	: data1 <= weights[3662];
				12'd3663	: data1 <= weights[3663];
				12'd3664	: data1 <= weights[3664];
				12'd3665	: data1 <= weights[3665];
				12'd3666	: data1 <= weights[3666];
				12'd3667	: data1 <= weights[3667];
				12'd3668	: data1 <= weights[3668];
				12'd3669	: data1 <= weights[3669];
				12'd3670	: data1 <= weights[3670];
				12'd3671	: data1 <= weights[3671];
				12'd3672	: data1 <= weights[3672];
				12'd3673	: data1 <= weights[3673];
				12'd3674	: data1 <= weights[3674];
				12'd3675	: data1 <= weights[3675];
				12'd3676	: data1 <= weights[3676];
				12'd3677	: data1 <= weights[3677];
				12'd3678	: data1 <= weights[3678];
				12'd3679	: data1 <= weights[3679];
				12'd3680	: data1 <= weights[3680];
				12'd3681	: data1 <= weights[3681];
				12'd3682	: data1 <= weights[3682];
				12'd3683	: data1 <= weights[3683];
				12'd3684	: data1 <= weights[3684];
				12'd3685	: data1 <= weights[3685];
				12'd3686	: data1 <= weights[3686];
				12'd3687	: data1 <= weights[3687];
				12'd3688	: data1 <= weights[3688];
				12'd3689	: data1 <= weights[3689];
				12'd3690	: data1 <= weights[3690];
				12'd3691	: data1 <= weights[3691];
				12'd3692	: data1 <= weights[3692];
				12'd3693	: data1 <= weights[3693];
				12'd3694	: data1 <= weights[3694];
				12'd3695	: data1 <= weights[3695];
				12'd3696	: data1 <= weights[3696];
				12'd3697	: data1 <= weights[3697];
				12'd3698	: data1 <= weights[3698];
				12'd3699	: data1 <= weights[3699];
				12'd3700	: data1 <= weights[3700];
				12'd3701	: data1 <= weights[3701];
				12'd3702	: data1 <= weights[3702];
				12'd3703	: data1 <= weights[3703];
				12'd3704	: data1 <= weights[3704];
				12'd3705	: data1 <= weights[3705];
				12'd3706	: data1 <= weights[3706];
				12'd3707	: data1 <= weights[3707];
				12'd3708	: data1 <= weights[3708];
				12'd3709	: data1 <= weights[3709];
				12'd3710	: data1 <= weights[3710];
				12'd3711	: data1 <= weights[3711];
				12'd3712	: data1 <= weights[3712];
				12'd3713	: data1 <= weights[3713];
				12'd3714	: data1 <= weights[3714];
				12'd3715	: data1 <= weights[3715];
				12'd3716	: data1 <= weights[3716];
				12'd3717	: data1 <= weights[3717];
				12'd3718	: data1 <= weights[3718];
				12'd3719	: data1 <= weights[3719];
				12'd3720	: data1 <= weights[3720];
				12'd3721	: data1 <= weights[3721];
				12'd3722	: data1 <= weights[3722];
				12'd3723	: data1 <= weights[3723];
				12'd3724	: data1 <= weights[3724];
				12'd3725	: data1 <= weights[3725];
				12'd3726	: data1 <= weights[3726];
				12'd3727	: data1 <= weights[3727];
				12'd3728	: data1 <= weights[3728];
				12'd3729	: data1 <= weights[3729];
				12'd3730	: data1 <= weights[3730];
				12'd3731	: data1 <= weights[3731];
				12'd3732	: data1 <= weights[3732];
				12'd3733	: data1 <= weights[3733];
				12'd3734	: data1 <= weights[3734];
				12'd3735	: data1 <= weights[3735];
				12'd3736	: data1 <= weights[3736];
				12'd3737	: data1 <= weights[3737];
				12'd3738	: data1 <= weights[3738];
				12'd3739	: data1 <= weights[3739];
				12'd3740	: data1 <= weights[3740];
				12'd3741	: data1 <= weights[3741];
				12'd3742	: data1 <= weights[3742];
				12'd3743	: data1 <= weights[3743];
				12'd3744	: data1 <= weights[3744];
				12'd3745	: data1 <= weights[3745];
				12'd3746	: data1 <= weights[3746];
				12'd3747	: data1 <= weights[3747];
				12'd3748	: data1 <= weights[3748];
				12'd3749	: data1 <= weights[3749];
				12'd3750	: data1 <= weights[3750];
				12'd3751	: data1 <= weights[3751];
				12'd3752	: data1 <= weights[3752];
				12'd3753	: data1 <= weights[3753];
				12'd3754	: data1 <= weights[3754];
				12'd3755	: data1 <= weights[3755];
				12'd3756	: data1 <= weights[3756];
				12'd3757	: data1 <= weights[3757];
				12'd3758	: data1 <= weights[3758];
				12'd3759	: data1 <= weights[3759];
				12'd3760	: data1 <= weights[3760];
				12'd3761	: data1 <= weights[3761];
				12'd3762	: data1 <= weights[3762];
				12'd3763	: data1 <= weights[3763];
				12'd3764	: data1 <= weights[3764];
				12'd3765	: data1 <= weights[3765];
				12'd3766	: data1 <= weights[3766];
				12'd3767	: data1 <= weights[3767];
				12'd3768	: data1 <= weights[3768];
				12'd3769	: data1 <= weights[3769];
				12'd3770	: data1 <= weights[3770];
				12'd3771	: data1 <= weights[3771];
				12'd3772	: data1 <= weights[3772];
				12'd3773	: data1 <= weights[3773];
				12'd3774	: data1 <= weights[3774];
				12'd3775	: data1 <= weights[3775];
				12'd3776	: data1 <= weights[3776];
				12'd3777	: data1 <= weights[3777];
				12'd3778	: data1 <= weights[3778];
				12'd3779	: data1 <= weights[3779];
				12'd3780	: data1 <= weights[3780];
				12'd3781	: data1 <= weights[3781];
				12'd3782	: data1 <= weights[3782];
				12'd3783	: data1 <= weights[3783];
				12'd3784	: data1 <= weights[3784];
				12'd3785	: data1 <= weights[3785];
				12'd3786	: data1 <= weights[3786];
				12'd3787	: data1 <= weights[3787];
				12'd3788	: data1 <= weights[3788];
				12'd3789	: data1 <= weights[3789];
				12'd3790	: data1 <= weights[3790];
				12'd3791	: data1 <= weights[3791];
				12'd3792	: data1 <= weights[3792];
				12'd3793	: data1 <= weights[3793];
				12'd3794	: data1 <= weights[3794];
				12'd3795	: data1 <= weights[3795];
				12'd3796	: data1 <= weights[3796];
				12'd3797	: data1 <= weights[3797];
				12'd3798	: data1 <= weights[3798];
				12'd3799	: data1 <= weights[3799];
				12'd3800	: data1 <= weights[3800];
				12'd3801	: data1 <= weights[3801];
				12'd3802	: data1 <= weights[3802];
				12'd3803	: data1 <= weights[3803];
				12'd3804	: data1 <= weights[3804];
				12'd3805	: data1 <= weights[3805];
				12'd3806	: data1 <= weights[3806];
				12'd3807	: data1 <= weights[3807];
				12'd3808	: data1 <= weights[3808];
				12'd3809	: data1 <= weights[3809];
				12'd3810	: data1 <= weights[3810];
				12'd3811	: data1 <= weights[3811];
				12'd3812	: data1 <= weights[3812];
				12'd3813	: data1 <= weights[3813];
				12'd3814	: data1 <= weights[3814];
				12'd3815	: data1 <= weights[3815];
				12'd3816	: data1 <= weights[3816];
				12'd3817	: data1 <= weights[3817];
				12'd3818	: data1 <= weights[3818];
				12'd3819	: data1 <= weights[3819];
				12'd3820	: data1 <= weights[3820];
				12'd3821	: data1 <= weights[3821];
				12'd3822	: data1 <= weights[3822];
				12'd3823	: data1 <= weights[3823];
				12'd3824	: data1 <= weights[3824];
				12'd3825	: data1 <= weights[3825];
				12'd3826	: data1 <= weights[3826];
				12'd3827	: data1 <= weights[3827];
				12'd3828	: data1 <= weights[3828];
				12'd3829	: data1 <= weights[3829];
				12'd3830	: data1 <= weights[3830];
				12'd3831	: data1 <= weights[3831];
				12'd3832	: data1 <= weights[3832];
				12'd3833	: data1 <= weights[3833];
				12'd3834	: data1 <= weights[3834];
				12'd3835	: data1 <= weights[3835];
				12'd3836	: data1 <= weights[3836];
				12'd3837	: data1 <= weights[3837];
				12'd3838	: data1 <= weights[3838];
				12'd3839	: data1 <= weights[3839];
				12'd3840	: data1 <= weights[3840];
				12'd3841	: data1 <= weights[3841];
				12'd3842	: data1 <= weights[3842];
				12'd3843	: data1 <= weights[3843];
				12'd3844	: data1 <= weights[3844];
				12'd3845	: data1 <= weights[3845];
				12'd3846	: data1 <= weights[3846];
				12'd3847	: data1 <= weights[3847];
				12'd3848	: data1 <= weights[3848];
				12'd3849	: data1 <= weights[3849];
				12'd3850	: data1 <= weights[3850];
				12'd3851	: data1 <= weights[3851];
				12'd3852	: data1 <= weights[3852];
				12'd3853	: data1 <= weights[3853];
				12'd3854	: data1 <= weights[3854];
				12'd3855	: data1 <= weights[3855];
				12'd3856	: data1 <= weights[3856];
				12'd3857	: data1 <= weights[3857];
				12'd3858	: data1 <= weights[3858];
				12'd3859	: data1 <= weights[3859];
				12'd3860	: data1 <= weights[3860];
				12'd3861	: data1 <= weights[3861];
				12'd3862	: data1 <= weights[3862];
				12'd3863	: data1 <= weights[3863];
				12'd3864	: data1 <= weights[3864];
				12'd3865	: data1 <= weights[3865];
				12'd3866	: data1 <= weights[3866];
				12'd3867	: data1 <= weights[3867];
				12'd3868	: data1 <= weights[3868];
				12'd3869	: data1 <= weights[3869];
				12'd3870	: data1 <= weights[3870];
				12'd3871	: data1 <= weights[3871];
				12'd3872	: data1 <= weights[3872];
				12'd3873	: data1 <= weights[3873];
				12'd3874	: data1 <= weights[3874];
				12'd3875	: data1 <= weights[3875];
				12'd3876	: data1 <= weights[3876];
				12'd3877	: data1 <= weights[3877];
				12'd3878	: data1 <= weights[3878];
				12'd3879	: data1 <= weights[3879];
				12'd3880	: data1 <= weights[3880];
				12'd3881	: data1 <= weights[3881];
				12'd3882	: data1 <= weights[3882];
				12'd3883	: data1 <= weights[3883];
				12'd3884	: data1 <= weights[3884];
				12'd3885	: data1 <= weights[3885];
				12'd3886	: data1 <= weights[3886];
				12'd3887	: data1 <= weights[3887];
				12'd3888	: data1 <= weights[3888];
				12'd3889	: data1 <= weights[3889];
				12'd3890	: data1 <= weights[3890];
				12'd3891	: data1 <= weights[3891];
				12'd3892	: data1 <= weights[3892];
				12'd3893	: data1 <= weights[3893];
				12'd3894	: data1 <= weights[3894];
				12'd3895	: data1 <= weights[3895];
				12'd3896	: data1 <= weights[3896];
				12'd3897	: data1 <= weights[3897];
				12'd3898	: data1 <= weights[3898];
				12'd3899	: data1 <= weights[3899];
				12'd3900	: data1 <= weights[3900];
				12'd3901	: data1 <= weights[3901];
				12'd3902	: data1 <= weights[3902];
				12'd3903	: data1 <= weights[3903];
				12'd3904	: data1 <= weights[3904];
				12'd3905	: data1 <= weights[3905];
				12'd3906	: data1 <= weights[3906];
				12'd3907	: data1 <= weights[3907];
				12'd3908	: data1 <= weights[3908];
				12'd3909	: data1 <= weights[3909];
				12'd3910	: data1 <= weights[3910];
				12'd3911	: data1 <= weights[3911];
				12'd3912	: data1 <= weights[3912];
				12'd3913	: data1 <= weights[3913];
				12'd3914	: data1 <= weights[3914];
				12'd3915	: data1 <= weights[3915];
				12'd3916	: data1 <= weights[3916];
				12'd3917	: data1 <= weights[3917];
				12'd3918	: data1 <= weights[3918];
				12'd3919	: data1 <= weights[3919];
				12'd3920	: data1 <= weights[3920];
				12'd3921	: data1 <= weights[3921];
				12'd3922	: data1 <= weights[3922];
				12'd3923	: data1 <= weights[3923];
				12'd3924	: data1 <= weights[3924];
				12'd3925	: data1 <= weights[3925];
				12'd3926	: data1 <= weights[3926];
				12'd3927	: data1 <= weights[3927];
				12'd3928	: data1 <= weights[3928];
				12'd3929	: data1 <= weights[3929];
				12'd3930	: data1 <= weights[3930];
				12'd3931	: data1 <= weights[3931];
				12'd3932	: data1 <= weights[3932];
				12'd3933	: data1 <= weights[3933];
				12'd3934	: data1 <= weights[3934];
				12'd3935	: data1 <= weights[3935];
				12'd3936	: data1 <= weights[3936];
				12'd3937	: data1 <= weights[3937];
				12'd3938	: data1 <= weights[3938];
				12'd3939	: data1 <= weights[3939];
				12'd3940	: data1 <= weights[3940];
				12'd3941	: data1 <= weights[3941];
				12'd3942	: data1 <= weights[3942];
				12'd3943	: data1 <= weights[3943];
				12'd3944	: data1 <= weights[3944];
				12'd3945	: data1 <= weights[3945];
				12'd3946	: data1 <= weights[3946];
				12'd3947	: data1 <= weights[3947];
				12'd3948	: data1 <= weights[3948];
				12'd3949	: data1 <= weights[3949];
				12'd3950	: data1 <= weights[3950];
				12'd3951	: data1 <= weights[3951];
				12'd3952	: data1 <= weights[3952];
				12'd3953	: data1 <= weights[3953];
				12'd3954	: data1 <= weights[3954];
				12'd3955	: data1 <= weights[3955];
				12'd3956	: data1 <= weights[3956];
				12'd3957	: data1 <= weights[3957];
				12'd3958	: data1 <= weights[3958];
				12'd3959	: data1 <= weights[3959];
				12'd3960	: data1 <= weights[3960];
				12'd3961	: data1 <= weights[3961];
				12'd3962	: data1 <= weights[3962];
				12'd3963	: data1 <= weights[3963];
				12'd3964	: data1 <= weights[3964];
				12'd3965	: data1 <= weights[3965];
				12'd3966	: data1 <= weights[3966];
				12'd3967	: data1 <= weights[3967];
				12'd3968	: data1 <= weights[3968];
				12'd3969	: data1 <= weights[3969];
				12'd3970	: data1 <= weights[3970];
				12'd3971	: data1 <= weights[3971];
				12'd3972	: data1 <= weights[3972];
				12'd3973	: data1 <= weights[3973];
				12'd3974	: data1 <= weights[3974];
				12'd3975	: data1 <= weights[3975];
				12'd3976	: data1 <= weights[3976];
				12'd3977	: data1 <= weights[3977];
				12'd3978	: data1 <= weights[3978];
				12'd3979	: data1 <= weights[3979];
				12'd3980	: data1 <= weights[3980];
				12'd3981	: data1 <= weights[3981];
				12'd3982	: data1 <= weights[3982];
				12'd3983	: data1 <= weights[3983];
				12'd3984	: data1 <= weights[3984];
				12'd3985	: data1 <= weights[3985];
				12'd3986	: data1 <= weights[3986];
				12'd3987	: data1 <= weights[3987];
				12'd3988	: data1 <= weights[3988];
				12'd3989	: data1 <= weights[3989];
				12'd3990	: data1 <= weights[3990];
				12'd3991	: data1 <= weights[3991];
				12'd3992	: data1 <= weights[3992];
				12'd3993	: data1 <= weights[3993];
				12'd3994	: data1 <= weights[3994];
				12'd3995	: data1 <= weights[3995];
				12'd3996	: data1 <= weights[3996];
				12'd3997	: data1 <= weights[3997];
				12'd3998	: data1 <= weights[3998];
				12'd3999	: data1 <= weights[3999];
				12'd4000	: data1 <= weights[4000];
				12'd4001	: data1 <= weights[4001];
				12'd4002	: data1 <= weights[4002];
				12'd4003	: data1 <= weights[4003];
				12'd4004	: data1 <= weights[4004];
				12'd4005	: data1 <= weights[4005];
				12'd4006	: data1 <= weights[4006];
				12'd4007	: data1 <= weights[4007];
				12'd4008	: data1 <= weights[4008];
				12'd4009	: data1 <= weights[4009];
				12'd4010	: data1 <= weights[4010];
				12'd4011	: data1 <= weights[4011];
				12'd4012	: data1 <= weights[4012];
				12'd4013	: data1 <= weights[4013];
				12'd4014	: data1 <= weights[4014];
				12'd4015	: data1 <= weights[4015];
				12'd4016	: data1 <= weights[4016];
				12'd4017	: data1 <= weights[4017];
				12'd4018	: data1 <= weights[4018];
				12'd4019	: data1 <= weights[4019];
				12'd4020	: data1 <= weights[4020];
				12'd4021	: data1 <= weights[4021];
				12'd4022	: data1 <= weights[4022];
				12'd4023	: data1 <= weights[4023];
				12'd4024	: data1 <= weights[4024];
				12'd4025	: data1 <= weights[4025];
				12'd4026	: data1 <= weights[4026];
				12'd4027	: data1 <= weights[4027];
				12'd4028	: data1 <= weights[4028];
				12'd4029	: data1 <= weights[4029];
				12'd4030	: data1 <= weights[4030];
				12'd4031	: data1 <= weights[4031];
				12'd4032	: data1 <= weights[4032];
				12'd4033	: data1 <= weights[4033];
				12'd4034	: data1 <= weights[4034];
				12'd4035	: data1 <= weights[4035];
				12'd4036	: data1 <= weights[4036];
				12'd4037	: data1 <= weights[4037];
				12'd4038	: data1 <= weights[4038];
				12'd4039	: data1 <= weights[4039];
				12'd4040	: data1 <= weights[4040];
				12'd4041	: data1 <= weights[4041];
				12'd4042	: data1 <= weights[4042];
				12'd4043	: data1 <= weights[4043];
				12'd4044	: data1 <= weights[4044];
				12'd4045	: data1 <= weights[4045];
				12'd4046	: data1 <= weights[4046];
				12'd4047	: data1 <= weights[4047];
				12'd4048	: data1 <= weights[4048];
				12'd4049	: data1 <= weights[4049];
				12'd4050	: data1 <= weights[4050];
				default		: data1 <= 16'd0;
			endcase
		end else begin
			data1 <= data1;
		end
	end


	always @(negedge(clk)) begin
		if(enable) begin
			case(address)
				12'd0		: data2 <= weights[1];
				12'd1		: data2 <= weights[2];
				12'd2		: data2 <= weights[3];
				12'd3		: data2 <= weights[4];
				12'd4		: data2 <= weights[5];
				12'd5		: data2 <= weights[6];
				12'd6		: data2 <= weights[7];
				12'd7		: data2 <= weights[8];
				12'd8		: data2 <= weights[9];
				12'd9		: data2 <= weights[10];
				12'd10		: data2 <= weights[11];
				12'd11		: data2 <= weights[12];
				12'd12		: data2 <= weights[13];
				12'd13		: data2 <= weights[14];
				12'd14		: data2 <= weights[15];
				12'd15		: data2 <= weights[16];
				12'd16		: data2 <= weights[17];
				12'd17		: data2 <= weights[18];
				12'd18		: data2 <= weights[19];
				12'd19		: data2 <= weights[20];
				12'd20		: data2 <= weights[21];
				12'd21		: data2 <= weights[22];
				12'd22		: data2 <= weights[23];
				12'd23		: data2 <= weights[24];
				12'd24		: data2 <= weights[25];
				12'd25		: data2 <= weights[26];
				12'd26		: data2 <= weights[27];
				12'd27		: data2 <= weights[28];
				12'd28		: data2 <= weights[29];
				12'd29		: data2 <= weights[30];
				12'd30		: data2 <= weights[31];
				12'd31		: data2 <= weights[32];
				12'd32		: data2 <= weights[33];
				12'd33		: data2 <= weights[34];
				12'd34		: data2 <= weights[35];
				12'd35		: data2 <= weights[36];
				12'd36		: data2 <= weights[37];
				12'd37		: data2 <= weights[38];
				12'd38		: data2 <= weights[39];
				12'd39		: data2 <= weights[40];
				12'd40		: data2 <= weights[41];
				12'd41		: data2 <= weights[42];
				12'd42		: data2 <= weights[43];
				12'd43		: data2 <= weights[44];
				12'd44		: data2 <= weights[45];
				12'd45		: data2 <= weights[46];
				12'd46		: data2 <= weights[47];
				12'd47		: data2 <= weights[48];
				12'd48		: data2 <= weights[49];
				12'd49		: data2 <= weights[50];
				12'd50		: data2 <= weights[51];
				12'd51		: data2 <= weights[52];
				12'd52		: data2 <= weights[53];
				12'd53		: data2 <= weights[54];
				12'd54		: data2 <= weights[55];
				12'd55		: data2 <= weights[56];
				12'd56		: data2 <= weights[57];
				12'd57		: data2 <= weights[58];
				12'd58		: data2 <= weights[59];
				12'd59		: data2 <= weights[60];
				12'd60		: data2 <= weights[61];
				12'd61		: data2 <= weights[62];
				12'd62		: data2 <= weights[63];
				12'd63		: data2 <= weights[64];
				12'd64		: data2 <= weights[65];
				12'd65		: data2 <= weights[66];
				12'd66		: data2 <= weights[67];
				12'd67		: data2 <= weights[68];
				12'd68		: data2 <= weights[69];
				12'd69		: data2 <= weights[70];
				12'd70		: data2 <= weights[71];
				12'd71		: data2 <= weights[72];
				12'd72		: data2 <= weights[73];
				12'd73		: data2 <= weights[74];
				12'd74		: data2 <= weights[75];
				12'd75		: data2 <= weights[76];
				12'd76		: data2 <= weights[77];
				12'd77		: data2 <= weights[78];
				12'd78		: data2 <= weights[79];
				12'd79		: data2 <= weights[80];
				12'd80		: data2 <= weights[81];
				12'd81		: data2 <= weights[82];
				12'd82		: data2 <= weights[83];
				12'd83		: data2 <= weights[84];
				12'd84		: data2 <= weights[85];
				12'd85		: data2 <= weights[86];
				12'd86		: data2 <= weights[87];
				12'd87		: data2 <= weights[88];
				12'd88		: data2 <= weights[89];
				12'd89		: data2 <= weights[90];
				12'd90		: data2 <= weights[91];
				12'd91		: data2 <= weights[92];
				12'd92		: data2 <= weights[93];
				12'd93		: data2 <= weights[94];
				12'd94		: data2 <= weights[95];
				12'd95		: data2 <= weights[96];
				12'd96		: data2 <= weights[97];
				12'd97		: data2 <= weights[98];
				12'd98		: data2 <= weights[99];
				12'd99		: data2 <= weights[100];
				12'd100		: data2 <= weights[101];
				12'd101		: data2 <= weights[102];
				12'd102		: data2 <= weights[103];
				12'd103		: data2 <= weights[104];
				12'd104		: data2 <= weights[105];
				12'd105		: data2 <= weights[106];
				12'd106		: data2 <= weights[107];
				12'd107		: data2 <= weights[108];
				12'd108		: data2 <= weights[109];
				12'd109		: data2 <= weights[110];
				12'd110		: data2 <= weights[111];
				12'd111		: data2 <= weights[112];
				12'd112		: data2 <= weights[113];
				12'd113		: data2 <= weights[114];
				12'd114		: data2 <= weights[115];
				12'd115		: data2 <= weights[116];
				12'd116		: data2 <= weights[117];
				12'd117		: data2 <= weights[118];
				12'd118		: data2 <= weights[119];
				12'd119		: data2 <= weights[120];
				12'd120		: data2 <= weights[121];
				12'd121		: data2 <= weights[122];
				12'd122		: data2 <= weights[123];
				12'd123		: data2 <= weights[124];
				12'd124		: data2 <= weights[125];
				12'd125		: data2 <= weights[126];
				12'd126		: data2 <= weights[127];
				12'd127		: data2 <= weights[128];
				12'd128		: data2 <= weights[129];
				12'd129		: data2 <= weights[130];
				12'd130		: data2 <= weights[131];
				12'd131		: data2 <= weights[132];
				12'd132		: data2 <= weights[133];
				12'd133		: data2 <= weights[134];
				12'd134		: data2 <= weights[135];
				12'd135		: data2 <= weights[136];
				12'd136		: data2 <= weights[137];
				12'd137		: data2 <= weights[138];
				12'd138		: data2 <= weights[139];
				12'd139		: data2 <= weights[140];
				12'd140		: data2 <= weights[141];
				12'd141		: data2 <= weights[142];
				12'd142		: data2 <= weights[143];
				12'd143		: data2 <= weights[144];
				12'd144		: data2 <= weights[145];
				12'd145		: data2 <= weights[146];
				12'd146		: data2 <= weights[147];
				12'd147		: data2 <= weights[148];
				12'd148		: data2 <= weights[149];
				12'd149		: data2 <= weights[150];
				12'd150		: data2 <= weights[151];
				12'd151		: data2 <= weights[152];
				12'd152		: data2 <= weights[153];
				12'd153		: data2 <= weights[154];
				12'd154		: data2 <= weights[155];
				12'd155		: data2 <= weights[156];
				12'd156		: data2 <= weights[157];
				12'd157		: data2 <= weights[158];
				12'd158		: data2 <= weights[159];
				12'd159		: data2 <= weights[160];
				12'd160		: data2 <= weights[161];
				12'd161		: data2 <= weights[162];
				12'd162		: data2 <= weights[163];
				12'd163		: data2 <= weights[164];
				12'd164		: data2 <= weights[165];
				12'd165		: data2 <= weights[166];
				12'd166		: data2 <= weights[167];
				12'd167		: data2 <= weights[168];
				12'd168		: data2 <= weights[169];
				12'd169		: data2 <= weights[170];
				12'd170		: data2 <= weights[171];
				12'd171		: data2 <= weights[172];
				12'd172		: data2 <= weights[173];
				12'd173		: data2 <= weights[174];
				12'd174		: data2 <= weights[175];
				12'd175		: data2 <= weights[176];
				12'd176		: data2 <= weights[177];
				12'd177		: data2 <= weights[178];
				12'd178		: data2 <= weights[179];
				12'd179		: data2 <= weights[180];
				12'd180		: data2 <= weights[181];
				12'd181		: data2 <= weights[182];
				12'd182		: data2 <= weights[183];
				12'd183		: data2 <= weights[184];
				12'd184		: data2 <= weights[185];
				12'd185		: data2 <= weights[186];
				12'd186		: data2 <= weights[187];
				12'd187		: data2 <= weights[188];
				12'd188		: data2 <= weights[189];
				12'd189		: data2 <= weights[190];
				12'd190		: data2 <= weights[191];
				12'd191		: data2 <= weights[192];
				12'd192		: data2 <= weights[193];
				12'd193		: data2 <= weights[194];
				12'd194		: data2 <= weights[195];
				12'd195		: data2 <= weights[196];
				12'd196		: data2 <= weights[197];
				12'd197		: data2 <= weights[198];
				12'd198		: data2 <= weights[199];
				12'd199		: data2 <= weights[200];
				12'd200		: data2 <= weights[201];
				12'd201		: data2 <= weights[202];
				12'd202		: data2 <= weights[203];
				12'd203		: data2 <= weights[204];
				12'd204		: data2 <= weights[205];
				12'd205		: data2 <= weights[206];
				12'd206		: data2 <= weights[207];
				12'd207		: data2 <= weights[208];
				12'd208		: data2 <= weights[209];
				12'd209		: data2 <= weights[210];
				12'd210		: data2 <= weights[211];
				12'd211		: data2 <= weights[212];
				12'd212		: data2 <= weights[213];
				12'd213		: data2 <= weights[214];
				12'd214		: data2 <= weights[215];
				12'd215		: data2 <= weights[216];
				12'd216		: data2 <= weights[217];
				12'd217		: data2 <= weights[218];
				12'd218		: data2 <= weights[219];
				12'd219		: data2 <= weights[220];
				12'd220		: data2 <= weights[221];
				12'd221		: data2 <= weights[222];
				12'd222		: data2 <= weights[223];
				12'd223		: data2 <= weights[224];
				12'd224		: data2 <= weights[225];
				12'd225		: data2 <= weights[226];
				12'd226		: data2 <= weights[227];
				12'd227		: data2 <= weights[228];
				12'd228		: data2 <= weights[229];
				12'd229		: data2 <= weights[230];
				12'd230		: data2 <= weights[231];
				12'd231		: data2 <= weights[232];
				12'd232		: data2 <= weights[233];
				12'd233		: data2 <= weights[234];
				12'd234		: data2 <= weights[235];
				12'd235		: data2 <= weights[236];
				12'd236		: data2 <= weights[237];
				12'd237		: data2 <= weights[238];
				12'd238		: data2 <= weights[239];
				12'd239		: data2 <= weights[240];
				12'd240		: data2 <= weights[241];
				12'd241		: data2 <= weights[242];
				12'd242		: data2 <= weights[243];
				12'd243		: data2 <= weights[244];
				12'd244		: data2 <= weights[245];
				12'd245		: data2 <= weights[246];
				12'd246		: data2 <= weights[247];
				12'd247		: data2 <= weights[248];
				12'd248		: data2 <= weights[249];
				12'd249		: data2 <= weights[250];
				12'd250		: data2 <= weights[251];
				12'd251		: data2 <= weights[252];
				12'd252		: data2 <= weights[253];
				12'd253		: data2 <= weights[254];
				12'd254		: data2 <= weights[255];
				12'd255		: data2 <= weights[256];
				12'd256		: data2 <= weights[257];
				12'd257		: data2 <= weights[258];
				12'd258		: data2 <= weights[259];
				12'd259		: data2 <= weights[260];
				12'd260		: data2 <= weights[261];
				12'd261		: data2 <= weights[262];
				12'd262		: data2 <= weights[263];
				12'd263		: data2 <= weights[264];
				12'd264		: data2 <= weights[265];
				12'd265		: data2 <= weights[266];
				12'd266		: data2 <= weights[267];
				12'd267		: data2 <= weights[268];
				12'd268		: data2 <= weights[269];
				12'd269		: data2 <= weights[270];
				12'd270		: data2 <= weights[271];
				12'd271		: data2 <= weights[272];
				12'd272		: data2 <= weights[273];
				12'd273		: data2 <= weights[274];
				12'd274		: data2 <= weights[275];
				12'd275		: data2 <= weights[276];
				12'd276		: data2 <= weights[277];
				12'd277		: data2 <= weights[278];
				12'd278		: data2 <= weights[279];
				12'd279		: data2 <= weights[280];
				12'd280		: data2 <= weights[281];
				12'd281		: data2 <= weights[282];
				12'd282		: data2 <= weights[283];
				12'd283		: data2 <= weights[284];
				12'd284		: data2 <= weights[285];
				12'd285		: data2 <= weights[286];
				12'd286		: data2 <= weights[287];
				12'd287		: data2 <= weights[288];
				12'd288		: data2 <= weights[289];
				12'd289		: data2 <= weights[290];
				12'd290		: data2 <= weights[291];
				12'd291		: data2 <= weights[292];
				12'd292		: data2 <= weights[293];
				12'd293		: data2 <= weights[294];
				12'd294		: data2 <= weights[295];
				12'd295		: data2 <= weights[296];
				12'd296		: data2 <= weights[297];
				12'd297		: data2 <= weights[298];
				12'd298		: data2 <= weights[299];
				12'd299		: data2 <= weights[300];
				12'd300		: data2 <= weights[301];
				12'd301		: data2 <= weights[302];
				12'd302		: data2 <= weights[303];
				12'd303		: data2 <= weights[304];
				12'd304		: data2 <= weights[305];
				12'd305		: data2 <= weights[306];
				12'd306		: data2 <= weights[307];
				12'd307		: data2 <= weights[308];
				12'd308		: data2 <= weights[309];
				12'd309		: data2 <= weights[310];
				12'd310		: data2 <= weights[311];
				12'd311		: data2 <= weights[312];
				12'd312		: data2 <= weights[313];
				12'd313		: data2 <= weights[314];
				12'd314		: data2 <= weights[315];
				12'd315		: data2 <= weights[316];
				12'd316		: data2 <= weights[317];
				12'd317		: data2 <= weights[318];
				12'd318		: data2 <= weights[319];
				12'd319		: data2 <= weights[320];
				12'd320		: data2 <= weights[321];
				12'd321		: data2 <= weights[322];
				12'd322		: data2 <= weights[323];
				12'd323		: data2 <= weights[324];
				12'd324		: data2 <= weights[325];
				12'd325		: data2 <= weights[326];
				12'd326		: data2 <= weights[327];
				12'd327		: data2 <= weights[328];
				12'd328		: data2 <= weights[329];
				12'd329		: data2 <= weights[330];
				12'd330		: data2 <= weights[331];
				12'd331		: data2 <= weights[332];
				12'd332		: data2 <= weights[333];
				12'd333		: data2 <= weights[334];
				12'd334		: data2 <= weights[335];
				12'd335		: data2 <= weights[336];
				12'd336		: data2 <= weights[337];
				12'd337		: data2 <= weights[338];
				12'd338		: data2 <= weights[339];
				12'd339		: data2 <= weights[340];
				12'd340		: data2 <= weights[341];
				12'd341		: data2 <= weights[342];
				12'd342		: data2 <= weights[343];
				12'd343		: data2 <= weights[344];
				12'd344		: data2 <= weights[345];
				12'd345		: data2 <= weights[346];
				12'd346		: data2 <= weights[347];
				12'd347		: data2 <= weights[348];
				12'd348		: data2 <= weights[349];
				12'd349		: data2 <= weights[350];
				12'd350		: data2 <= weights[351];
				12'd351		: data2 <= weights[352];
				12'd352		: data2 <= weights[353];
				12'd353		: data2 <= weights[354];
				12'd354		: data2 <= weights[355];
				12'd355		: data2 <= weights[356];
				12'd356		: data2 <= weights[357];
				12'd357		: data2 <= weights[358];
				12'd358		: data2 <= weights[359];
				12'd359		: data2 <= weights[360];
				12'd360		: data2 <= weights[361];
				12'd361		: data2 <= weights[362];
				12'd362		: data2 <= weights[363];
				12'd363		: data2 <= weights[364];
				12'd364		: data2 <= weights[365];
				12'd365		: data2 <= weights[366];
				12'd366		: data2 <= weights[367];
				12'd367		: data2 <= weights[368];
				12'd368		: data2 <= weights[369];
				12'd369		: data2 <= weights[370];
				12'd370		: data2 <= weights[371];
				12'd371		: data2 <= weights[372];
				12'd372		: data2 <= weights[373];
				12'd373		: data2 <= weights[374];
				12'd374		: data2 <= weights[375];
				12'd375		: data2 <= weights[376];
				12'd376		: data2 <= weights[377];
				12'd377		: data2 <= weights[378];
				12'd378		: data2 <= weights[379];
				12'd379		: data2 <= weights[380];
				12'd380		: data2 <= weights[381];
				12'd381		: data2 <= weights[382];
				12'd382		: data2 <= weights[383];
				12'd383		: data2 <= weights[384];
				12'd384		: data2 <= weights[385];
				12'd385		: data2 <= weights[386];
				12'd386		: data2 <= weights[387];
				12'd387		: data2 <= weights[388];
				12'd388		: data2 <= weights[389];
				12'd389		: data2 <= weights[390];
				12'd390		: data2 <= weights[391];
				12'd391		: data2 <= weights[392];
				12'd392		: data2 <= weights[393];
				12'd393		: data2 <= weights[394];
				12'd394		: data2 <= weights[395];
				12'd395		: data2 <= weights[396];
				12'd396		: data2 <= weights[397];
				12'd397		: data2 <= weights[398];
				12'd398		: data2 <= weights[399];
				12'd399		: data2 <= weights[400];
				12'd400		: data2 <= weights[401];
				12'd401		: data2 <= weights[402];
				12'd402		: data2 <= weights[403];
				12'd403		: data2 <= weights[404];
				12'd404		: data2 <= weights[405];
				12'd405		: data2 <= weights[406];
				12'd406		: data2 <= weights[407];
				12'd407		: data2 <= weights[408];
				12'd408		: data2 <= weights[409];
				12'd409		: data2 <= weights[410];
				12'd410		: data2 <= weights[411];
				12'd411		: data2 <= weights[412];
				12'd412		: data2 <= weights[413];
				12'd413		: data2 <= weights[414];
				12'd414		: data2 <= weights[415];
				12'd415		: data2 <= weights[416];
				12'd416		: data2 <= weights[417];
				12'd417		: data2 <= weights[418];
				12'd418		: data2 <= weights[419];
				12'd419		: data2 <= weights[420];
				12'd420		: data2 <= weights[421];
				12'd421		: data2 <= weights[422];
				12'd422		: data2 <= weights[423];
				12'd423		: data2 <= weights[424];
				12'd424		: data2 <= weights[425];
				12'd425		: data2 <= weights[426];
				12'd426		: data2 <= weights[427];
				12'd427		: data2 <= weights[428];
				12'd428		: data2 <= weights[429];
				12'd429		: data2 <= weights[430];
				12'd430		: data2 <= weights[431];
				12'd431		: data2 <= weights[432];
				12'd432		: data2 <= weights[433];
				12'd433		: data2 <= weights[434];
				12'd434		: data2 <= weights[435];
				12'd435		: data2 <= weights[436];
				12'd436		: data2 <= weights[437];
				12'd437		: data2 <= weights[438];
				12'd438		: data2 <= weights[439];
				12'd439		: data2 <= weights[440];
				12'd440		: data2 <= weights[441];
				12'd441		: data2 <= weights[442];
				12'd442		: data2 <= weights[443];
				12'd443		: data2 <= weights[444];
				12'd444		: data2 <= weights[445];
				12'd445		: data2 <= weights[446];
				12'd446		: data2 <= weights[447];
				12'd447		: data2 <= weights[448];
				12'd448		: data2 <= weights[449];
				12'd449		: data2 <= weights[450];
				12'd450		: data2 <= weights[451];
				12'd451		: data2 <= weights[452];
				12'd452		: data2 <= weights[453];
				12'd453		: data2 <= weights[454];
				12'd454		: data2 <= weights[455];
				12'd455		: data2 <= weights[456];
				12'd456		: data2 <= weights[457];
				12'd457		: data2 <= weights[458];
				12'd458		: data2 <= weights[459];
				12'd459		: data2 <= weights[460];
				12'd460		: data2 <= weights[461];
				12'd461		: data2 <= weights[462];
				12'd462		: data2 <= weights[463];
				12'd463		: data2 <= weights[464];
				12'd464		: data2 <= weights[465];
				12'd465		: data2 <= weights[466];
				12'd466		: data2 <= weights[467];
				12'd467		: data2 <= weights[468];
				12'd468		: data2 <= weights[469];
				12'd469		: data2 <= weights[470];
				12'd470		: data2 <= weights[471];
				12'd471		: data2 <= weights[472];
				12'd472		: data2 <= weights[473];
				12'd473		: data2 <= weights[474];
				12'd474		: data2 <= weights[475];
				12'd475		: data2 <= weights[476];
				12'd476		: data2 <= weights[477];
				12'd477		: data2 <= weights[478];
				12'd478		: data2 <= weights[479];
				12'd479		: data2 <= weights[480];
				12'd480		: data2 <= weights[481];
				12'd481		: data2 <= weights[482];
				12'd482		: data2 <= weights[483];
				12'd483		: data2 <= weights[484];
				12'd484		: data2 <= weights[485];
				12'd485		: data2 <= weights[486];
				12'd486		: data2 <= weights[487];
				12'd487		: data2 <= weights[488];
				12'd488		: data2 <= weights[489];
				12'd489		: data2 <= weights[490];
				12'd490		: data2 <= weights[491];
				12'd491		: data2 <= weights[492];
				12'd492		: data2 <= weights[493];
				12'd493		: data2 <= weights[494];
				12'd494		: data2 <= weights[495];
				12'd495		: data2 <= weights[496];
				12'd496		: data2 <= weights[497];
				12'd497		: data2 <= weights[498];
				12'd498		: data2 <= weights[499];
				12'd499		: data2 <= weights[500];
				12'd500		: data2 <= weights[501];
				12'd501		: data2 <= weights[502];
				12'd502		: data2 <= weights[503];
				12'd503		: data2 <= weights[504];
				12'd504		: data2 <= weights[505];
				12'd505		: data2 <= weights[506];
				12'd506		: data2 <= weights[507];
				12'd507		: data2 <= weights[508];
				12'd508		: data2 <= weights[509];
				12'd509		: data2 <= weights[510];
				12'd510		: data2 <= weights[511];
				12'd511		: data2 <= weights[512];
				12'd512		: data2 <= weights[513];
				12'd513		: data2 <= weights[514];
				12'd514		: data2 <= weights[515];
				12'd515		: data2 <= weights[516];
				12'd516		: data2 <= weights[517];
				12'd517		: data2 <= weights[518];
				12'd518		: data2 <= weights[519];
				12'd519		: data2 <= weights[520];
				12'd520		: data2 <= weights[521];
				12'd521		: data2 <= weights[522];
				12'd522		: data2 <= weights[523];
				12'd523		: data2 <= weights[524];
				12'd524		: data2 <= weights[525];
				12'd525		: data2 <= weights[526];
				12'd526		: data2 <= weights[527];
				12'd527		: data2 <= weights[528];
				12'd528		: data2 <= weights[529];
				12'd529		: data2 <= weights[530];
				12'd530		: data2 <= weights[531];
				12'd531		: data2 <= weights[532];
				12'd532		: data2 <= weights[533];
				12'd533		: data2 <= weights[534];
				12'd534		: data2 <= weights[535];
				12'd535		: data2 <= weights[536];
				12'd536		: data2 <= weights[537];
				12'd537		: data2 <= weights[538];
				12'd538		: data2 <= weights[539];
				12'd539		: data2 <= weights[540];
				12'd540		: data2 <= weights[541];
				12'd541		: data2 <= weights[542];
				12'd542		: data2 <= weights[543];
				12'd543		: data2 <= weights[544];
				12'd544		: data2 <= weights[545];
				12'd545		: data2 <= weights[546];
				12'd546		: data2 <= weights[547];
				12'd547		: data2 <= weights[548];
				12'd548		: data2 <= weights[549];
				12'd549		: data2 <= weights[550];
				12'd550		: data2 <= weights[551];
				12'd551		: data2 <= weights[552];
				12'd552		: data2 <= weights[553];
				12'd553		: data2 <= weights[554];
				12'd554		: data2 <= weights[555];
				12'd555		: data2 <= weights[556];
				12'd556		: data2 <= weights[557];
				12'd557		: data2 <= weights[558];
				12'd558		: data2 <= weights[559];
				12'd559		: data2 <= weights[560];
				12'd560		: data2 <= weights[561];
				12'd561		: data2 <= weights[562];
				12'd562		: data2 <= weights[563];
				12'd563		: data2 <= weights[564];
				12'd564		: data2 <= weights[565];
				12'd565		: data2 <= weights[566];
				12'd566		: data2 <= weights[567];
				12'd567		: data2 <= weights[568];
				12'd568		: data2 <= weights[569];
				12'd569		: data2 <= weights[570];
				12'd570		: data2 <= weights[571];
				12'd571		: data2 <= weights[572];
				12'd572		: data2 <= weights[573];
				12'd573		: data2 <= weights[574];
				12'd574		: data2 <= weights[575];
				12'd575		: data2 <= weights[576];
				12'd576		: data2 <= weights[577];
				12'd577		: data2 <= weights[578];
				12'd578		: data2 <= weights[579];
				12'd579		: data2 <= weights[580];
				12'd580		: data2 <= weights[581];
				12'd581		: data2 <= weights[582];
				12'd582		: data2 <= weights[583];
				12'd583		: data2 <= weights[584];
				12'd584		: data2 <= weights[585];
				12'd585		: data2 <= weights[586];
				12'd586		: data2 <= weights[587];
				12'd587		: data2 <= weights[588];
				12'd588		: data2 <= weights[589];
				12'd589		: data2 <= weights[590];
				12'd590		: data2 <= weights[591];
				12'd591		: data2 <= weights[592];
				12'd592		: data2 <= weights[593];
				12'd593		: data2 <= weights[594];
				12'd594		: data2 <= weights[595];
				12'd595		: data2 <= weights[596];
				12'd596		: data2 <= weights[597];
				12'd597		: data2 <= weights[598];
				12'd598		: data2 <= weights[599];
				12'd599		: data2 <= weights[600];
				12'd600		: data2 <= weights[601];
				12'd601		: data2 <= weights[602];
				12'd602		: data2 <= weights[603];
				12'd603		: data2 <= weights[604];
				12'd604		: data2 <= weights[605];
				12'd605		: data2 <= weights[606];
				12'd606		: data2 <= weights[607];
				12'd607		: data2 <= weights[608];
				12'd608		: data2 <= weights[609];
				12'd609		: data2 <= weights[610];
				12'd610		: data2 <= weights[611];
				12'd611		: data2 <= weights[612];
				12'd612		: data2 <= weights[613];
				12'd613		: data2 <= weights[614];
				12'd614		: data2 <= weights[615];
				12'd615		: data2 <= weights[616];
				12'd616		: data2 <= weights[617];
				12'd617		: data2 <= weights[618];
				12'd618		: data2 <= weights[619];
				12'd619		: data2 <= weights[620];
				12'd620		: data2 <= weights[621];
				12'd621		: data2 <= weights[622];
				12'd622		: data2 <= weights[623];
				12'd623		: data2 <= weights[624];
				12'd624		: data2 <= weights[625];
				12'd625		: data2 <= weights[626];
				12'd626		: data2 <= weights[627];
				12'd627		: data2 <= weights[628];
				12'd628		: data2 <= weights[629];
				12'd629		: data2 <= weights[630];
				12'd630		: data2 <= weights[631];
				12'd631		: data2 <= weights[632];
				12'd632		: data2 <= weights[633];
				12'd633		: data2 <= weights[634];
				12'd634		: data2 <= weights[635];
				12'd635		: data2 <= weights[636];
				12'd636		: data2 <= weights[637];
				12'd637		: data2 <= weights[638];
				12'd638		: data2 <= weights[639];
				12'd639		: data2 <= weights[640];
				12'd640		: data2 <= weights[641];
				12'd641		: data2 <= weights[642];
				12'd642		: data2 <= weights[643];
				12'd643		: data2 <= weights[644];
				12'd644		: data2 <= weights[645];
				12'd645		: data2 <= weights[646];
				12'd646		: data2 <= weights[647];
				12'd647		: data2 <= weights[648];
				12'd648		: data2 <= weights[649];
				12'd649		: data2 <= weights[650];
				12'd650		: data2 <= weights[651];
				12'd651		: data2 <= weights[652];
				12'd652		: data2 <= weights[653];
				12'd653		: data2 <= weights[654];
				12'd654		: data2 <= weights[655];
				12'd655		: data2 <= weights[656];
				12'd656		: data2 <= weights[657];
				12'd657		: data2 <= weights[658];
				12'd658		: data2 <= weights[659];
				12'd659		: data2 <= weights[660];
				12'd660		: data2 <= weights[661];
				12'd661		: data2 <= weights[662];
				12'd662		: data2 <= weights[663];
				12'd663		: data2 <= weights[664];
				12'd664		: data2 <= weights[665];
				12'd665		: data2 <= weights[666];
				12'd666		: data2 <= weights[667];
				12'd667		: data2 <= weights[668];
				12'd668		: data2 <= weights[669];
				12'd669		: data2 <= weights[670];
				12'd670		: data2 <= weights[671];
				12'd671		: data2 <= weights[672];
				12'd672		: data2 <= weights[673];
				12'd673		: data2 <= weights[674];
				12'd674		: data2 <= weights[675];
				12'd675		: data2 <= weights[676];
				12'd676		: data2 <= weights[677];
				12'd677		: data2 <= weights[678];
				12'd678		: data2 <= weights[679];
				12'd679		: data2 <= weights[680];
				12'd680		: data2 <= weights[681];
				12'd681		: data2 <= weights[682];
				12'd682		: data2 <= weights[683];
				12'd683		: data2 <= weights[684];
				12'd684		: data2 <= weights[685];
				12'd685		: data2 <= weights[686];
				12'd686		: data2 <= weights[687];
				12'd687		: data2 <= weights[688];
				12'd688		: data2 <= weights[689];
				12'd689		: data2 <= weights[690];
				12'd690		: data2 <= weights[691];
				12'd691		: data2 <= weights[692];
				12'd692		: data2 <= weights[693];
				12'd693		: data2 <= weights[694];
				12'd694		: data2 <= weights[695];
				12'd695		: data2 <= weights[696];
				12'd696		: data2 <= weights[697];
				12'd697		: data2 <= weights[698];
				12'd698		: data2 <= weights[699];
				12'd699		: data2 <= weights[700];
				12'd700		: data2 <= weights[701];
				12'd701		: data2 <= weights[702];
				12'd702		: data2 <= weights[703];
				12'd703		: data2 <= weights[704];
				12'd704		: data2 <= weights[705];
				12'd705		: data2 <= weights[706];
				12'd706		: data2 <= weights[707];
				12'd707		: data2 <= weights[708];
				12'd708		: data2 <= weights[709];
				12'd709		: data2 <= weights[710];
				12'd710		: data2 <= weights[711];
				12'd711		: data2 <= weights[712];
				12'd712		: data2 <= weights[713];
				12'd713		: data2 <= weights[714];
				12'd714		: data2 <= weights[715];
				12'd715		: data2 <= weights[716];
				12'd716		: data2 <= weights[717];
				12'd717		: data2 <= weights[718];
				12'd718		: data2 <= weights[719];
				12'd719		: data2 <= weights[720];
				12'd720		: data2 <= weights[721];
				12'd721		: data2 <= weights[722];
				12'd722		: data2 <= weights[723];
				12'd723		: data2 <= weights[724];
				12'd724		: data2 <= weights[725];
				12'd725		: data2 <= weights[726];
				12'd726		: data2 <= weights[727];
				12'd727		: data2 <= weights[728];
				12'd728		: data2 <= weights[729];
				12'd729		: data2 <= weights[730];
				12'd730		: data2 <= weights[731];
				12'd731		: data2 <= weights[732];
				12'd732		: data2 <= weights[733];
				12'd733		: data2 <= weights[734];
				12'd734		: data2 <= weights[735];
				12'd735		: data2 <= weights[736];
				12'd736		: data2 <= weights[737];
				12'd737		: data2 <= weights[738];
				12'd738		: data2 <= weights[739];
				12'd739		: data2 <= weights[740];
				12'd740		: data2 <= weights[741];
				12'd741		: data2 <= weights[742];
				12'd742		: data2 <= weights[743];
				12'd743		: data2 <= weights[744];
				12'd744		: data2 <= weights[745];
				12'd745		: data2 <= weights[746];
				12'd746		: data2 <= weights[747];
				12'd747		: data2 <= weights[748];
				12'd748		: data2 <= weights[749];
				12'd749		: data2 <= weights[750];
				12'd750		: data2 <= weights[751];
				12'd751		: data2 <= weights[752];
				12'd752		: data2 <= weights[753];
				12'd753		: data2 <= weights[754];
				12'd754		: data2 <= weights[755];
				12'd755		: data2 <= weights[756];
				12'd756		: data2 <= weights[757];
				12'd757		: data2 <= weights[758];
				12'd758		: data2 <= weights[759];
				12'd759		: data2 <= weights[760];
				12'd760		: data2 <= weights[761];
				12'd761		: data2 <= weights[762];
				12'd762		: data2 <= weights[763];
				12'd763		: data2 <= weights[764];
				12'd764		: data2 <= weights[765];
				12'd765		: data2 <= weights[766];
				12'd766		: data2 <= weights[767];
				12'd767		: data2 <= weights[768];
				12'd768		: data2 <= weights[769];
				12'd769		: data2 <= weights[770];
				12'd770		: data2 <= weights[771];
				12'd771		: data2 <= weights[772];
				12'd772		: data2 <= weights[773];
				12'd773		: data2 <= weights[774];
				12'd774		: data2 <= weights[775];
				12'd775		: data2 <= weights[776];
				12'd776		: data2 <= weights[777];
				12'd777		: data2 <= weights[778];
				12'd778		: data2 <= weights[779];
				12'd779		: data2 <= weights[780];
				12'd780		: data2 <= weights[781];
				12'd781		: data2 <= weights[782];
				12'd782		: data2 <= weights[783];
				12'd783		: data2 <= weights[784];
				12'd784		: data2 <= weights[785];
				12'd785		: data2 <= weights[786];
				12'd786		: data2 <= weights[787];
				12'd787		: data2 <= weights[788];
				12'd788		: data2 <= weights[789];
				12'd789		: data2 <= weights[790];
				12'd790		: data2 <= weights[791];
				12'd791		: data2 <= weights[792];
				12'd792		: data2 <= weights[793];
				12'd793		: data2 <= weights[794];
				12'd794		: data2 <= weights[795];
				12'd795		: data2 <= weights[796];
				12'd796		: data2 <= weights[797];
				12'd797		: data2 <= weights[798];
				12'd798		: data2 <= weights[799];
				12'd799		: data2 <= weights[800];
				12'd800		: data2 <= weights[801];
				12'd801		: data2 <= weights[802];
				12'd802		: data2 <= weights[803];
				12'd803		: data2 <= weights[804];
				12'd804		: data2 <= weights[805];
				12'd805		: data2 <= weights[806];
				12'd806		: data2 <= weights[807];
				12'd807		: data2 <= weights[808];
				12'd808		: data2 <= weights[809];
				12'd809		: data2 <= weights[810];
				12'd810		: data2 <= weights[811];
				12'd811		: data2 <= weights[812];
				12'd812		: data2 <= weights[813];
				12'd813		: data2 <= weights[814];
				12'd814		: data2 <= weights[815];
				12'd815		: data2 <= weights[816];
				12'd816		: data2 <= weights[817];
				12'd817		: data2 <= weights[818];
				12'd818		: data2 <= weights[819];
				12'd819		: data2 <= weights[820];
				12'd820		: data2 <= weights[821];
				12'd821		: data2 <= weights[822];
				12'd822		: data2 <= weights[823];
				12'd823		: data2 <= weights[824];
				12'd824		: data2 <= weights[825];
				12'd825		: data2 <= weights[826];
				12'd826		: data2 <= weights[827];
				12'd827		: data2 <= weights[828];
				12'd828		: data2 <= weights[829];
				12'd829		: data2 <= weights[830];
				12'd830		: data2 <= weights[831];
				12'd831		: data2 <= weights[832];
				12'd832		: data2 <= weights[833];
				12'd833		: data2 <= weights[834];
				12'd834		: data2 <= weights[835];
				12'd835		: data2 <= weights[836];
				12'd836		: data2 <= weights[837];
				12'd837		: data2 <= weights[838];
				12'd838		: data2 <= weights[839];
				12'd839		: data2 <= weights[840];
				12'd840		: data2 <= weights[841];
				12'd841		: data2 <= weights[842];
				12'd842		: data2 <= weights[843];
				12'd843		: data2 <= weights[844];
				12'd844		: data2 <= weights[845];
				12'd845		: data2 <= weights[846];
				12'd846		: data2 <= weights[847];
				12'd847		: data2 <= weights[848];
				12'd848		: data2 <= weights[849];
				12'd849		: data2 <= weights[850];
				12'd850		: data2 <= weights[851];
				12'd851		: data2 <= weights[852];
				12'd852		: data2 <= weights[853];
				12'd853		: data2 <= weights[854];
				12'd854		: data2 <= weights[855];
				12'd855		: data2 <= weights[856];
				12'd856		: data2 <= weights[857];
				12'd857		: data2 <= weights[858];
				12'd858		: data2 <= weights[859];
				12'd859		: data2 <= weights[860];
				12'd860		: data2 <= weights[861];
				12'd861		: data2 <= weights[862];
				12'd862		: data2 <= weights[863];
				12'd863		: data2 <= weights[864];
				12'd864		: data2 <= weights[865];
				12'd865		: data2 <= weights[866];
				12'd866		: data2 <= weights[867];
				12'd867		: data2 <= weights[868];
				12'd868		: data2 <= weights[869];
				12'd869		: data2 <= weights[870];
				12'd870		: data2 <= weights[871];
				12'd871		: data2 <= weights[872];
				12'd872		: data2 <= weights[873];
				12'd873		: data2 <= weights[874];
				12'd874		: data2 <= weights[875];
				12'd875		: data2 <= weights[876];
				12'd876		: data2 <= weights[877];
				12'd877		: data2 <= weights[878];
				12'd878		: data2 <= weights[879];
				12'd879		: data2 <= weights[880];
				12'd880		: data2 <= weights[881];
				12'd881		: data2 <= weights[882];
				12'd882		: data2 <= weights[883];
				12'd883		: data2 <= weights[884];
				12'd884		: data2 <= weights[885];
				12'd885		: data2 <= weights[886];
				12'd886		: data2 <= weights[887];
				12'd887		: data2 <= weights[888];
				12'd888		: data2 <= weights[889];
				12'd889		: data2 <= weights[890];
				12'd890		: data2 <= weights[891];
				12'd891		: data2 <= weights[892];
				12'd892		: data2 <= weights[893];
				12'd893		: data2 <= weights[894];
				12'd894		: data2 <= weights[895];
				12'd895		: data2 <= weights[896];
				12'd896		: data2 <= weights[897];
				12'd897		: data2 <= weights[898];
				12'd898		: data2 <= weights[899];
				12'd899		: data2 <= weights[900];
				12'd900		: data2 <= weights[901];
				12'd901		: data2 <= weights[902];
				12'd902		: data2 <= weights[903];
				12'd903		: data2 <= weights[904];
				12'd904		: data2 <= weights[905];
				12'd905		: data2 <= weights[906];
				12'd906		: data2 <= weights[907];
				12'd907		: data2 <= weights[908];
				12'd908		: data2 <= weights[909];
				12'd909		: data2 <= weights[910];
				12'd910		: data2 <= weights[911];
				12'd911		: data2 <= weights[912];
				12'd912		: data2 <= weights[913];
				12'd913		: data2 <= weights[914];
				12'd914		: data2 <= weights[915];
				12'd915		: data2 <= weights[916];
				12'd916		: data2 <= weights[917];
				12'd917		: data2 <= weights[918];
				12'd918		: data2 <= weights[919];
				12'd919		: data2 <= weights[920];
				12'd920		: data2 <= weights[921];
				12'd921		: data2 <= weights[922];
				12'd922		: data2 <= weights[923];
				12'd923		: data2 <= weights[924];
				12'd924		: data2 <= weights[925];
				12'd925		: data2 <= weights[926];
				12'd926		: data2 <= weights[927];
				12'd927		: data2 <= weights[928];
				12'd928		: data2 <= weights[929];
				12'd929		: data2 <= weights[930];
				12'd930		: data2 <= weights[931];
				12'd931		: data2 <= weights[932];
				12'd932		: data2 <= weights[933];
				12'd933		: data2 <= weights[934];
				12'd934		: data2 <= weights[935];
				12'd935		: data2 <= weights[936];
				12'd936		: data2 <= weights[937];
				12'd937		: data2 <= weights[938];
				12'd938		: data2 <= weights[939];
				12'd939		: data2 <= weights[940];
				12'd940		: data2 <= weights[941];
				12'd941		: data2 <= weights[942];
				12'd942		: data2 <= weights[943];
				12'd943		: data2 <= weights[944];
				12'd944		: data2 <= weights[945];
				12'd945		: data2 <= weights[946];
				12'd946		: data2 <= weights[947];
				12'd947		: data2 <= weights[948];
				12'd948		: data2 <= weights[949];
				12'd949		: data2 <= weights[950];
				12'd950		: data2 <= weights[951];
				12'd951		: data2 <= weights[952];
				12'd952		: data2 <= weights[953];
				12'd953		: data2 <= weights[954];
				12'd954		: data2 <= weights[955];
				12'd955		: data2 <= weights[956];
				12'd956		: data2 <= weights[957];
				12'd957		: data2 <= weights[958];
				12'd958		: data2 <= weights[959];
				12'd959		: data2 <= weights[960];
				12'd960		: data2 <= weights[961];
				12'd961		: data2 <= weights[962];
				12'd962		: data2 <= weights[963];
				12'd963		: data2 <= weights[964];
				12'd964		: data2 <= weights[965];
				12'd965		: data2 <= weights[966];
				12'd966		: data2 <= weights[967];
				12'd967		: data2 <= weights[968];
				12'd968		: data2 <= weights[969];
				12'd969		: data2 <= weights[970];
				12'd970		: data2 <= weights[971];
				12'd971		: data2 <= weights[972];
				12'd972		: data2 <= weights[973];
				12'd973		: data2 <= weights[974];
				12'd974		: data2 <= weights[975];
				12'd975		: data2 <= weights[976];
				12'd976		: data2 <= weights[977];
				12'd977		: data2 <= weights[978];
				12'd978		: data2 <= weights[979];
				12'd979		: data2 <= weights[980];
				12'd980		: data2 <= weights[981];
				12'd981		: data2 <= weights[982];
				12'd982		: data2 <= weights[983];
				12'd983		: data2 <= weights[984];
				12'd984		: data2 <= weights[985];
				12'd985		: data2 <= weights[986];
				12'd986		: data2 <= weights[987];
				12'd987		: data2 <= weights[988];
				12'd988		: data2 <= weights[989];
				12'd989		: data2 <= weights[990];
				12'd990		: data2 <= weights[991];
				12'd991		: data2 <= weights[992];
				12'd992		: data2 <= weights[993];
				12'd993		: data2 <= weights[994];
				12'd994		: data2 <= weights[995];
				12'd995		: data2 <= weights[996];
				12'd996		: data2 <= weights[997];
				12'd997		: data2 <= weights[998];
				12'd998		: data2 <= weights[999];
				12'd999		: data2 <= weights[1000];
				12'd1000	: data2 <= weights[1001];
				12'd1001	: data2 <= weights[1002];
				12'd1002	: data2 <= weights[1003];
				12'd1003	: data2 <= weights[1004];
				12'd1004	: data2 <= weights[1005];
				12'd1005	: data2 <= weights[1006];
				12'd1006	: data2 <= weights[1007];
				12'd1007	: data2 <= weights[1008];
				12'd1008	: data2 <= weights[1009];
				12'd1009	: data2 <= weights[1010];
				12'd1010	: data2 <= weights[1011];
				12'd1011	: data2 <= weights[1012];
				12'd1012	: data2 <= weights[1013];
				12'd1013	: data2 <= weights[1014];
				12'd1014	: data2 <= weights[1015];
				12'd1015	: data2 <= weights[1016];
				12'd1016	: data2 <= weights[1017];
				12'd1017	: data2 <= weights[1018];
				12'd1018	: data2 <= weights[1019];
				12'd1019	: data2 <= weights[1020];
				12'd1020	: data2 <= weights[1021];
				12'd1021	: data2 <= weights[1022];
				12'd1022	: data2 <= weights[1023];
				12'd1023	: data2 <= weights[1024];
				12'd1024	: data2 <= weights[1025];
				12'd1025	: data2 <= weights[1026];
				12'd1026	: data2 <= weights[1027];
				12'd1027	: data2 <= weights[1028];
				12'd1028	: data2 <= weights[1029];
				12'd1029	: data2 <= weights[1030];
				12'd1030	: data2 <= weights[1031];
				12'd1031	: data2 <= weights[1032];
				12'd1032	: data2 <= weights[1033];
				12'd1033	: data2 <= weights[1034];
				12'd1034	: data2 <= weights[1035];
				12'd1035	: data2 <= weights[1036];
				12'd1036	: data2 <= weights[1037];
				12'd1037	: data2 <= weights[1038];
				12'd1038	: data2 <= weights[1039];
				12'd1039	: data2 <= weights[1040];
				12'd1040	: data2 <= weights[1041];
				12'd1041	: data2 <= weights[1042];
				12'd1042	: data2 <= weights[1043];
				12'd1043	: data2 <= weights[1044];
				12'd1044	: data2 <= weights[1045];
				12'd1045	: data2 <= weights[1046];
				12'd1046	: data2 <= weights[1047];
				12'd1047	: data2 <= weights[1048];
				12'd1048	: data2 <= weights[1049];
				12'd1049	: data2 <= weights[1050];
				12'd1050	: data2 <= weights[1051];
				12'd1051	: data2 <= weights[1052];
				12'd1052	: data2 <= weights[1053];
				12'd1053	: data2 <= weights[1054];
				12'd1054	: data2 <= weights[1055];
				12'd1055	: data2 <= weights[1056];
				12'd1056	: data2 <= weights[1057];
				12'd1057	: data2 <= weights[1058];
				12'd1058	: data2 <= weights[1059];
				12'd1059	: data2 <= weights[1060];
				12'd1060	: data2 <= weights[1061];
				12'd1061	: data2 <= weights[1062];
				12'd1062	: data2 <= weights[1063];
				12'd1063	: data2 <= weights[1064];
				12'd1064	: data2 <= weights[1065];
				12'd1065	: data2 <= weights[1066];
				12'd1066	: data2 <= weights[1067];
				12'd1067	: data2 <= weights[1068];
				12'd1068	: data2 <= weights[1069];
				12'd1069	: data2 <= weights[1070];
				12'd1070	: data2 <= weights[1071];
				12'd1071	: data2 <= weights[1072];
				12'd1072	: data2 <= weights[1073];
				12'd1073	: data2 <= weights[1074];
				12'd1074	: data2 <= weights[1075];
				12'd1075	: data2 <= weights[1076];
				12'd1076	: data2 <= weights[1077];
				12'd1077	: data2 <= weights[1078];
				12'd1078	: data2 <= weights[1079];
				12'd1079	: data2 <= weights[1080];
				12'd1080	: data2 <= weights[1081];
				12'd1081	: data2 <= weights[1082];
				12'd1082	: data2 <= weights[1083];
				12'd1083	: data2 <= weights[1084];
				12'd1084	: data2 <= weights[1085];
				12'd1085	: data2 <= weights[1086];
				12'd1086	: data2 <= weights[1087];
				12'd1087	: data2 <= weights[1088];
				12'd1088	: data2 <= weights[1089];
				12'd1089	: data2 <= weights[1090];
				12'd1090	: data2 <= weights[1091];
				12'd1091	: data2 <= weights[1092];
				12'd1092	: data2 <= weights[1093];
				12'd1093	: data2 <= weights[1094];
				12'd1094	: data2 <= weights[1095];
				12'd1095	: data2 <= weights[1096];
				12'd1096	: data2 <= weights[1097];
				12'd1097	: data2 <= weights[1098];
				12'd1098	: data2 <= weights[1099];
				12'd1099	: data2 <= weights[1100];
				12'd1100	: data2 <= weights[1101];
				12'd1101	: data2 <= weights[1102];
				12'd1102	: data2 <= weights[1103];
				12'd1103	: data2 <= weights[1104];
				12'd1104	: data2 <= weights[1105];
				12'd1105	: data2 <= weights[1106];
				12'd1106	: data2 <= weights[1107];
				12'd1107	: data2 <= weights[1108];
				12'd1108	: data2 <= weights[1109];
				12'd1109	: data2 <= weights[1110];
				12'd1110	: data2 <= weights[1111];
				12'd1111	: data2 <= weights[1112];
				12'd1112	: data2 <= weights[1113];
				12'd1113	: data2 <= weights[1114];
				12'd1114	: data2 <= weights[1115];
				12'd1115	: data2 <= weights[1116];
				12'd1116	: data2 <= weights[1117];
				12'd1117	: data2 <= weights[1118];
				12'd1118	: data2 <= weights[1119];
				12'd1119	: data2 <= weights[1120];
				12'd1120	: data2 <= weights[1121];
				12'd1121	: data2 <= weights[1122];
				12'd1122	: data2 <= weights[1123];
				12'd1123	: data2 <= weights[1124];
				12'd1124	: data2 <= weights[1125];
				12'd1125	: data2 <= weights[1126];
				12'd1126	: data2 <= weights[1127];
				12'd1127	: data2 <= weights[1128];
				12'd1128	: data2 <= weights[1129];
				12'd1129	: data2 <= weights[1130];
				12'd1130	: data2 <= weights[1131];
				12'd1131	: data2 <= weights[1132];
				12'd1132	: data2 <= weights[1133];
				12'd1133	: data2 <= weights[1134];
				12'd1134	: data2 <= weights[1135];
				12'd1135	: data2 <= weights[1136];
				12'd1136	: data2 <= weights[1137];
				12'd1137	: data2 <= weights[1138];
				12'd1138	: data2 <= weights[1139];
				12'd1139	: data2 <= weights[1140];
				12'd1140	: data2 <= weights[1141];
				12'd1141	: data2 <= weights[1142];
				12'd1142	: data2 <= weights[1143];
				12'd1143	: data2 <= weights[1144];
				12'd1144	: data2 <= weights[1145];
				12'd1145	: data2 <= weights[1146];
				12'd1146	: data2 <= weights[1147];
				12'd1147	: data2 <= weights[1148];
				12'd1148	: data2 <= weights[1149];
				12'd1149	: data2 <= weights[1150];
				12'd1150	: data2 <= weights[1151];
				12'd1151	: data2 <= weights[1152];
				12'd1152	: data2 <= weights[1153];
				12'd1153	: data2 <= weights[1154];
				12'd1154	: data2 <= weights[1155];
				12'd1155	: data2 <= weights[1156];
				12'd1156	: data2 <= weights[1157];
				12'd1157	: data2 <= weights[1158];
				12'd1158	: data2 <= weights[1159];
				12'd1159	: data2 <= weights[1160];
				12'd1160	: data2 <= weights[1161];
				12'd1161	: data2 <= weights[1162];
				12'd1162	: data2 <= weights[1163];
				12'd1163	: data2 <= weights[1164];
				12'd1164	: data2 <= weights[1165];
				12'd1165	: data2 <= weights[1166];
				12'd1166	: data2 <= weights[1167];
				12'd1167	: data2 <= weights[1168];
				12'd1168	: data2 <= weights[1169];
				12'd1169	: data2 <= weights[1170];
				12'd1170	: data2 <= weights[1171];
				12'd1171	: data2 <= weights[1172];
				12'd1172	: data2 <= weights[1173];
				12'd1173	: data2 <= weights[1174];
				12'd1174	: data2 <= weights[1175];
				12'd1175	: data2 <= weights[1176];
				12'd1176	: data2 <= weights[1177];
				12'd1177	: data2 <= weights[1178];
				12'd1178	: data2 <= weights[1179];
				12'd1179	: data2 <= weights[1180];
				12'd1180	: data2 <= weights[1181];
				12'd1181	: data2 <= weights[1182];
				12'd1182	: data2 <= weights[1183];
				12'd1183	: data2 <= weights[1184];
				12'd1184	: data2 <= weights[1185];
				12'd1185	: data2 <= weights[1186];
				12'd1186	: data2 <= weights[1187];
				12'd1187	: data2 <= weights[1188];
				12'd1188	: data2 <= weights[1189];
				12'd1189	: data2 <= weights[1190];
				12'd1190	: data2 <= weights[1191];
				12'd1191	: data2 <= weights[1192];
				12'd1192	: data2 <= weights[1193];
				12'd1193	: data2 <= weights[1194];
				12'd1194	: data2 <= weights[1195];
				12'd1195	: data2 <= weights[1196];
				12'd1196	: data2 <= weights[1197];
				12'd1197	: data2 <= weights[1198];
				12'd1198	: data2 <= weights[1199];
				12'd1199	: data2 <= weights[1200];
				12'd1200	: data2 <= weights[1201];
				12'd1201	: data2 <= weights[1202];
				12'd1202	: data2 <= weights[1203];
				12'd1203	: data2 <= weights[1204];
				12'd1204	: data2 <= weights[1205];
				12'd1205	: data2 <= weights[1206];
				12'd1206	: data2 <= weights[1207];
				12'd1207	: data2 <= weights[1208];
				12'd1208	: data2 <= weights[1209];
				12'd1209	: data2 <= weights[1210];
				12'd1210	: data2 <= weights[1211];
				12'd1211	: data2 <= weights[1212];
				12'd1212	: data2 <= weights[1213];
				12'd1213	: data2 <= weights[1214];
				12'd1214	: data2 <= weights[1215];
				12'd1215	: data2 <= weights[1216];
				12'd1216	: data2 <= weights[1217];
				12'd1217	: data2 <= weights[1218];
				12'd1218	: data2 <= weights[1219];
				12'd1219	: data2 <= weights[1220];
				12'd1220	: data2 <= weights[1221];
				12'd1221	: data2 <= weights[1222];
				12'd1222	: data2 <= weights[1223];
				12'd1223	: data2 <= weights[1224];
				12'd1224	: data2 <= weights[1225];
				12'd1225	: data2 <= weights[1226];
				12'd1226	: data2 <= weights[1227];
				12'd1227	: data2 <= weights[1228];
				12'd1228	: data2 <= weights[1229];
				12'd1229	: data2 <= weights[1230];
				12'd1230	: data2 <= weights[1231];
				12'd1231	: data2 <= weights[1232];
				12'd1232	: data2 <= weights[1233];
				12'd1233	: data2 <= weights[1234];
				12'd1234	: data2 <= weights[1235];
				12'd1235	: data2 <= weights[1236];
				12'd1236	: data2 <= weights[1237];
				12'd1237	: data2 <= weights[1238];
				12'd1238	: data2 <= weights[1239];
				12'd1239	: data2 <= weights[1240];
				12'd1240	: data2 <= weights[1241];
				12'd1241	: data2 <= weights[1242];
				12'd1242	: data2 <= weights[1243];
				12'd1243	: data2 <= weights[1244];
				12'd1244	: data2 <= weights[1245];
				12'd1245	: data2 <= weights[1246];
				12'd1246	: data2 <= weights[1247];
				12'd1247	: data2 <= weights[1248];
				12'd1248	: data2 <= weights[1249];
				12'd1249	: data2 <= weights[1250];
				12'd1250	: data2 <= weights[1251];
				12'd1251	: data2 <= weights[1252];
				12'd1252	: data2 <= weights[1253];
				12'd1253	: data2 <= weights[1254];
				12'd1254	: data2 <= weights[1255];
				12'd1255	: data2 <= weights[1256];
				12'd1256	: data2 <= weights[1257];
				12'd1257	: data2 <= weights[1258];
				12'd1258	: data2 <= weights[1259];
				12'd1259	: data2 <= weights[1260];
				12'd1260	: data2 <= weights[1261];
				12'd1261	: data2 <= weights[1262];
				12'd1262	: data2 <= weights[1263];
				12'd1263	: data2 <= weights[1264];
				12'd1264	: data2 <= weights[1265];
				12'd1265	: data2 <= weights[1266];
				12'd1266	: data2 <= weights[1267];
				12'd1267	: data2 <= weights[1268];
				12'd1268	: data2 <= weights[1269];
				12'd1269	: data2 <= weights[1270];
				12'd1270	: data2 <= weights[1271];
				12'd1271	: data2 <= weights[1272];
				12'd1272	: data2 <= weights[1273];
				12'd1273	: data2 <= weights[1274];
				12'd1274	: data2 <= weights[1275];
				12'd1275	: data2 <= weights[1276];
				12'd1276	: data2 <= weights[1277];
				12'd1277	: data2 <= weights[1278];
				12'd1278	: data2 <= weights[1279];
				12'd1279	: data2 <= weights[1280];
				12'd1280	: data2 <= weights[1281];
				12'd1281	: data2 <= weights[1282];
				12'd1282	: data2 <= weights[1283];
				12'd1283	: data2 <= weights[1284];
				12'd1284	: data2 <= weights[1285];
				12'd1285	: data2 <= weights[1286];
				12'd1286	: data2 <= weights[1287];
				12'd1287	: data2 <= weights[1288];
				12'd1288	: data2 <= weights[1289];
				12'd1289	: data2 <= weights[1290];
				12'd1290	: data2 <= weights[1291];
				12'd1291	: data2 <= weights[1292];
				12'd1292	: data2 <= weights[1293];
				12'd1293	: data2 <= weights[1294];
				12'd1294	: data2 <= weights[1295];
				12'd1295	: data2 <= weights[1296];
				12'd1296	: data2 <= weights[1297];
				12'd1297	: data2 <= weights[1298];
				12'd1298	: data2 <= weights[1299];
				12'd1299	: data2 <= weights[1300];
				12'd1300	: data2 <= weights[1301];
				12'd1301	: data2 <= weights[1302];
				12'd1302	: data2 <= weights[1303];
				12'd1303	: data2 <= weights[1304];
				12'd1304	: data2 <= weights[1305];
				12'd1305	: data2 <= weights[1306];
				12'd1306	: data2 <= weights[1307];
				12'd1307	: data2 <= weights[1308];
				12'd1308	: data2 <= weights[1309];
				12'd1309	: data2 <= weights[1310];
				12'd1310	: data2 <= weights[1311];
				12'd1311	: data2 <= weights[1312];
				12'd1312	: data2 <= weights[1313];
				12'd1313	: data2 <= weights[1314];
				12'd1314	: data2 <= weights[1315];
				12'd1315	: data2 <= weights[1316];
				12'd1316	: data2 <= weights[1317];
				12'd1317	: data2 <= weights[1318];
				12'd1318	: data2 <= weights[1319];
				12'd1319	: data2 <= weights[1320];
				12'd1320	: data2 <= weights[1321];
				12'd1321	: data2 <= weights[1322];
				12'd1322	: data2 <= weights[1323];
				12'd1323	: data2 <= weights[1324];
				12'd1324	: data2 <= weights[1325];
				12'd1325	: data2 <= weights[1326];
				12'd1326	: data2 <= weights[1327];
				12'd1327	: data2 <= weights[1328];
				12'd1328	: data2 <= weights[1329];
				12'd1329	: data2 <= weights[1330];
				12'd1330	: data2 <= weights[1331];
				12'd1331	: data2 <= weights[1332];
				12'd1332	: data2 <= weights[1333];
				12'd1333	: data2 <= weights[1334];
				12'd1334	: data2 <= weights[1335];
				12'd1335	: data2 <= weights[1336];
				12'd1336	: data2 <= weights[1337];
				12'd1337	: data2 <= weights[1338];
				12'd1338	: data2 <= weights[1339];
				12'd1339	: data2 <= weights[1340];
				12'd1340	: data2 <= weights[1341];
				12'd1341	: data2 <= weights[1342];
				12'd1342	: data2 <= weights[1343];
				12'd1343	: data2 <= weights[1344];
				12'd1344	: data2 <= weights[1345];
				12'd1345	: data2 <= weights[1346];
				12'd1346	: data2 <= weights[1347];
				12'd1347	: data2 <= weights[1348];
				12'd1348	: data2 <= weights[1349];
				12'd1349	: data2 <= weights[1350];
				12'd1350	: data2 <= weights[1351];
				12'd1351	: data2 <= weights[1352];
				12'd1352	: data2 <= weights[1353];
				12'd1353	: data2 <= weights[1354];
				12'd1354	: data2 <= weights[1355];
				12'd1355	: data2 <= weights[1356];
				12'd1356	: data2 <= weights[1357];
				12'd1357	: data2 <= weights[1358];
				12'd1358	: data2 <= weights[1359];
				12'd1359	: data2 <= weights[1360];
				12'd1360	: data2 <= weights[1361];
				12'd1361	: data2 <= weights[1362];
				12'd1362	: data2 <= weights[1363];
				12'd1363	: data2 <= weights[1364];
				12'd1364	: data2 <= weights[1365];
				12'd1365	: data2 <= weights[1366];
				12'd1366	: data2 <= weights[1367];
				12'd1367	: data2 <= weights[1368];
				12'd1368	: data2 <= weights[1369];
				12'd1369	: data2 <= weights[1370];
				12'd1370	: data2 <= weights[1371];
				12'd1371	: data2 <= weights[1372];
				12'd1372	: data2 <= weights[1373];
				12'd1373	: data2 <= weights[1374];
				12'd1374	: data2 <= weights[1375];
				12'd1375	: data2 <= weights[1376];
				12'd1376	: data2 <= weights[1377];
				12'd1377	: data2 <= weights[1378];
				12'd1378	: data2 <= weights[1379];
				12'd1379	: data2 <= weights[1380];
				12'd1380	: data2 <= weights[1381];
				12'd1381	: data2 <= weights[1382];
				12'd1382	: data2 <= weights[1383];
				12'd1383	: data2 <= weights[1384];
				12'd1384	: data2 <= weights[1385];
				12'd1385	: data2 <= weights[1386];
				12'd1386	: data2 <= weights[1387];
				12'd1387	: data2 <= weights[1388];
				12'd1388	: data2 <= weights[1389];
				12'd1389	: data2 <= weights[1390];
				12'd1390	: data2 <= weights[1391];
				12'd1391	: data2 <= weights[1392];
				12'd1392	: data2 <= weights[1393];
				12'd1393	: data2 <= weights[1394];
				12'd1394	: data2 <= weights[1395];
				12'd1395	: data2 <= weights[1396];
				12'd1396	: data2 <= weights[1397];
				12'd1397	: data2 <= weights[1398];
				12'd1398	: data2 <= weights[1399];
				12'd1399	: data2 <= weights[1400];
				12'd1400	: data2 <= weights[1401];
				12'd1401	: data2 <= weights[1402];
				12'd1402	: data2 <= weights[1403];
				12'd1403	: data2 <= weights[1404];
				12'd1404	: data2 <= weights[1405];
				12'd1405	: data2 <= weights[1406];
				12'd1406	: data2 <= weights[1407];
				12'd1407	: data2 <= weights[1408];
				12'd1408	: data2 <= weights[1409];
				12'd1409	: data2 <= weights[1410];
				12'd1410	: data2 <= weights[1411];
				12'd1411	: data2 <= weights[1412];
				12'd1412	: data2 <= weights[1413];
				12'd1413	: data2 <= weights[1414];
				12'd1414	: data2 <= weights[1415];
				12'd1415	: data2 <= weights[1416];
				12'd1416	: data2 <= weights[1417];
				12'd1417	: data2 <= weights[1418];
				12'd1418	: data2 <= weights[1419];
				12'd1419	: data2 <= weights[1420];
				12'd1420	: data2 <= weights[1421];
				12'd1421	: data2 <= weights[1422];
				12'd1422	: data2 <= weights[1423];
				12'd1423	: data2 <= weights[1424];
				12'd1424	: data2 <= weights[1425];
				12'd1425	: data2 <= weights[1426];
				12'd1426	: data2 <= weights[1427];
				12'd1427	: data2 <= weights[1428];
				12'd1428	: data2 <= weights[1429];
				12'd1429	: data2 <= weights[1430];
				12'd1430	: data2 <= weights[1431];
				12'd1431	: data2 <= weights[1432];
				12'd1432	: data2 <= weights[1433];
				12'd1433	: data2 <= weights[1434];
				12'd1434	: data2 <= weights[1435];
				12'd1435	: data2 <= weights[1436];
				12'd1436	: data2 <= weights[1437];
				12'd1437	: data2 <= weights[1438];
				12'd1438	: data2 <= weights[1439];
				12'd1439	: data2 <= weights[1440];
				12'd1440	: data2 <= weights[1441];
				12'd1441	: data2 <= weights[1442];
				12'd1442	: data2 <= weights[1443];
				12'd1443	: data2 <= weights[1444];
				12'd1444	: data2 <= weights[1445];
				12'd1445	: data2 <= weights[1446];
				12'd1446	: data2 <= weights[1447];
				12'd1447	: data2 <= weights[1448];
				12'd1448	: data2 <= weights[1449];
				12'd1449	: data2 <= weights[1450];
				12'd1450	: data2 <= weights[1451];
				12'd1451	: data2 <= weights[1452];
				12'd1452	: data2 <= weights[1453];
				12'd1453	: data2 <= weights[1454];
				12'd1454	: data2 <= weights[1455];
				12'd1455	: data2 <= weights[1456];
				12'd1456	: data2 <= weights[1457];
				12'd1457	: data2 <= weights[1458];
				12'd1458	: data2 <= weights[1459];
				12'd1459	: data2 <= weights[1460];
				12'd1460	: data2 <= weights[1461];
				12'd1461	: data2 <= weights[1462];
				12'd1462	: data2 <= weights[1463];
				12'd1463	: data2 <= weights[1464];
				12'd1464	: data2 <= weights[1465];
				12'd1465	: data2 <= weights[1466];
				12'd1466	: data2 <= weights[1467];
				12'd1467	: data2 <= weights[1468];
				12'd1468	: data2 <= weights[1469];
				12'd1469	: data2 <= weights[1470];
				12'd1470	: data2 <= weights[1471];
				12'd1471	: data2 <= weights[1472];
				12'd1472	: data2 <= weights[1473];
				12'd1473	: data2 <= weights[1474];
				12'd1474	: data2 <= weights[1475];
				12'd1475	: data2 <= weights[1476];
				12'd1476	: data2 <= weights[1477];
				12'd1477	: data2 <= weights[1478];
				12'd1478	: data2 <= weights[1479];
				12'd1479	: data2 <= weights[1480];
				12'd1480	: data2 <= weights[1481];
				12'd1481	: data2 <= weights[1482];
				12'd1482	: data2 <= weights[1483];
				12'd1483	: data2 <= weights[1484];
				12'd1484	: data2 <= weights[1485];
				12'd1485	: data2 <= weights[1486];
				12'd1486	: data2 <= weights[1487];
				12'd1487	: data2 <= weights[1488];
				12'd1488	: data2 <= weights[1489];
				12'd1489	: data2 <= weights[1490];
				12'd1490	: data2 <= weights[1491];
				12'd1491	: data2 <= weights[1492];
				12'd1492	: data2 <= weights[1493];
				12'd1493	: data2 <= weights[1494];
				12'd1494	: data2 <= weights[1495];
				12'd1495	: data2 <= weights[1496];
				12'd1496	: data2 <= weights[1497];
				12'd1497	: data2 <= weights[1498];
				12'd1498	: data2 <= weights[1499];
				12'd1499	: data2 <= weights[1500];
				12'd1500	: data2 <= weights[1501];
				12'd1501	: data2 <= weights[1502];
				12'd1502	: data2 <= weights[1503];
				12'd1503	: data2 <= weights[1504];
				12'd1504	: data2 <= weights[1505];
				12'd1505	: data2 <= weights[1506];
				12'd1506	: data2 <= weights[1507];
				12'd1507	: data2 <= weights[1508];
				12'd1508	: data2 <= weights[1509];
				12'd1509	: data2 <= weights[1510];
				12'd1510	: data2 <= weights[1511];
				12'd1511	: data2 <= weights[1512];
				12'd1512	: data2 <= weights[1513];
				12'd1513	: data2 <= weights[1514];
				12'd1514	: data2 <= weights[1515];
				12'd1515	: data2 <= weights[1516];
				12'd1516	: data2 <= weights[1517];
				12'd1517	: data2 <= weights[1518];
				12'd1518	: data2 <= weights[1519];
				12'd1519	: data2 <= weights[1520];
				12'd1520	: data2 <= weights[1521];
				12'd1521	: data2 <= weights[1522];
				12'd1522	: data2 <= weights[1523];
				12'd1523	: data2 <= weights[1524];
				12'd1524	: data2 <= weights[1525];
				12'd1525	: data2 <= weights[1526];
				12'd1526	: data2 <= weights[1527];
				12'd1527	: data2 <= weights[1528];
				12'd1528	: data2 <= weights[1529];
				12'd1529	: data2 <= weights[1530];
				12'd1530	: data2 <= weights[1531];
				12'd1531	: data2 <= weights[1532];
				12'd1532	: data2 <= weights[1533];
				12'd1533	: data2 <= weights[1534];
				12'd1534	: data2 <= weights[1535];
				12'd1535	: data2 <= weights[1536];
				12'd1536	: data2 <= weights[1537];
				12'd1537	: data2 <= weights[1538];
				12'd1538	: data2 <= weights[1539];
				12'd1539	: data2 <= weights[1540];
				12'd1540	: data2 <= weights[1541];
				12'd1541	: data2 <= weights[1542];
				12'd1542	: data2 <= weights[1543];
				12'd1543	: data2 <= weights[1544];
				12'd1544	: data2 <= weights[1545];
				12'd1545	: data2 <= weights[1546];
				12'd1546	: data2 <= weights[1547];
				12'd1547	: data2 <= weights[1548];
				12'd1548	: data2 <= weights[1549];
				12'd1549	: data2 <= weights[1550];
				12'd1550	: data2 <= weights[1551];
				12'd1551	: data2 <= weights[1552];
				12'd1552	: data2 <= weights[1553];
				12'd1553	: data2 <= weights[1554];
				12'd1554	: data2 <= weights[1555];
				12'd1555	: data2 <= weights[1556];
				12'd1556	: data2 <= weights[1557];
				12'd1557	: data2 <= weights[1558];
				12'd1558	: data2 <= weights[1559];
				12'd1559	: data2 <= weights[1560];
				12'd1560	: data2 <= weights[1561];
				12'd1561	: data2 <= weights[1562];
				12'd1562	: data2 <= weights[1563];
				12'd1563	: data2 <= weights[1564];
				12'd1564	: data2 <= weights[1565];
				12'd1565	: data2 <= weights[1566];
				12'd1566	: data2 <= weights[1567];
				12'd1567	: data2 <= weights[1568];
				12'd1568	: data2 <= weights[1569];
				12'd1569	: data2 <= weights[1570];
				12'd1570	: data2 <= weights[1571];
				12'd1571	: data2 <= weights[1572];
				12'd1572	: data2 <= weights[1573];
				12'd1573	: data2 <= weights[1574];
				12'd1574	: data2 <= weights[1575];
				12'd1575	: data2 <= weights[1576];
				12'd1576	: data2 <= weights[1577];
				12'd1577	: data2 <= weights[1578];
				12'd1578	: data2 <= weights[1579];
				12'd1579	: data2 <= weights[1580];
				12'd1580	: data2 <= weights[1581];
				12'd1581	: data2 <= weights[1582];
				12'd1582	: data2 <= weights[1583];
				12'd1583	: data2 <= weights[1584];
				12'd1584	: data2 <= weights[1585];
				12'd1585	: data2 <= weights[1586];
				12'd1586	: data2 <= weights[1587];
				12'd1587	: data2 <= weights[1588];
				12'd1588	: data2 <= weights[1589];
				12'd1589	: data2 <= weights[1590];
				12'd1590	: data2 <= weights[1591];
				12'd1591	: data2 <= weights[1592];
				12'd1592	: data2 <= weights[1593];
				12'd1593	: data2 <= weights[1594];
				12'd1594	: data2 <= weights[1595];
				12'd1595	: data2 <= weights[1596];
				12'd1596	: data2 <= weights[1597];
				12'd1597	: data2 <= weights[1598];
				12'd1598	: data2 <= weights[1599];
				12'd1599	: data2 <= weights[1600];
				12'd1600	: data2 <= weights[1601];
				12'd1601	: data2 <= weights[1602];
				12'd1602	: data2 <= weights[1603];
				12'd1603	: data2 <= weights[1604];
				12'd1604	: data2 <= weights[1605];
				12'd1605	: data2 <= weights[1606];
				12'd1606	: data2 <= weights[1607];
				12'd1607	: data2 <= weights[1608];
				12'd1608	: data2 <= weights[1609];
				12'd1609	: data2 <= weights[1610];
				12'd1610	: data2 <= weights[1611];
				12'd1611	: data2 <= weights[1612];
				12'd1612	: data2 <= weights[1613];
				12'd1613	: data2 <= weights[1614];
				12'd1614	: data2 <= weights[1615];
				12'd1615	: data2 <= weights[1616];
				12'd1616	: data2 <= weights[1617];
				12'd1617	: data2 <= weights[1618];
				12'd1618	: data2 <= weights[1619];
				12'd1619	: data2 <= weights[1620];
				12'd1620	: data2 <= weights[1621];
				12'd1621	: data2 <= weights[1622];
				12'd1622	: data2 <= weights[1623];
				12'd1623	: data2 <= weights[1624];
				12'd1624	: data2 <= weights[1625];
				12'd1625	: data2 <= weights[1626];
				12'd1626	: data2 <= weights[1627];
				12'd1627	: data2 <= weights[1628];
				12'd1628	: data2 <= weights[1629];
				12'd1629	: data2 <= weights[1630];
				12'd1630	: data2 <= weights[1631];
				12'd1631	: data2 <= weights[1632];
				12'd1632	: data2 <= weights[1633];
				12'd1633	: data2 <= weights[1634];
				12'd1634	: data2 <= weights[1635];
				12'd1635	: data2 <= weights[1636];
				12'd1636	: data2 <= weights[1637];
				12'd1637	: data2 <= weights[1638];
				12'd1638	: data2 <= weights[1639];
				12'd1639	: data2 <= weights[1640];
				12'd1640	: data2 <= weights[1641];
				12'd1641	: data2 <= weights[1642];
				12'd1642	: data2 <= weights[1643];
				12'd1643	: data2 <= weights[1644];
				12'd1644	: data2 <= weights[1645];
				12'd1645	: data2 <= weights[1646];
				12'd1646	: data2 <= weights[1647];
				12'd1647	: data2 <= weights[1648];
				12'd1648	: data2 <= weights[1649];
				12'd1649	: data2 <= weights[1650];
				12'd1650	: data2 <= weights[1651];
				12'd1651	: data2 <= weights[1652];
				12'd1652	: data2 <= weights[1653];
				12'd1653	: data2 <= weights[1654];
				12'd1654	: data2 <= weights[1655];
				12'd1655	: data2 <= weights[1656];
				12'd1656	: data2 <= weights[1657];
				12'd1657	: data2 <= weights[1658];
				12'd1658	: data2 <= weights[1659];
				12'd1659	: data2 <= weights[1660];
				12'd1660	: data2 <= weights[1661];
				12'd1661	: data2 <= weights[1662];
				12'd1662	: data2 <= weights[1663];
				12'd1663	: data2 <= weights[1664];
				12'd1664	: data2 <= weights[1665];
				12'd1665	: data2 <= weights[1666];
				12'd1666	: data2 <= weights[1667];
				12'd1667	: data2 <= weights[1668];
				12'd1668	: data2 <= weights[1669];
				12'd1669	: data2 <= weights[1670];
				12'd1670	: data2 <= weights[1671];
				12'd1671	: data2 <= weights[1672];
				12'd1672	: data2 <= weights[1673];
				12'd1673	: data2 <= weights[1674];
				12'd1674	: data2 <= weights[1675];
				12'd1675	: data2 <= weights[1676];
				12'd1676	: data2 <= weights[1677];
				12'd1677	: data2 <= weights[1678];
				12'd1678	: data2 <= weights[1679];
				12'd1679	: data2 <= weights[1680];
				12'd1680	: data2 <= weights[1681];
				12'd1681	: data2 <= weights[1682];
				12'd1682	: data2 <= weights[1683];
				12'd1683	: data2 <= weights[1684];
				12'd1684	: data2 <= weights[1685];
				12'd1685	: data2 <= weights[1686];
				12'd1686	: data2 <= weights[1687];
				12'd1687	: data2 <= weights[1688];
				12'd1688	: data2 <= weights[1689];
				12'd1689	: data2 <= weights[1690];
				12'd1690	: data2 <= weights[1691];
				12'd1691	: data2 <= weights[1692];
				12'd1692	: data2 <= weights[1693];
				12'd1693	: data2 <= weights[1694];
				12'd1694	: data2 <= weights[1695];
				12'd1695	: data2 <= weights[1696];
				12'd1696	: data2 <= weights[1697];
				12'd1697	: data2 <= weights[1698];
				12'd1698	: data2 <= weights[1699];
				12'd1699	: data2 <= weights[1700];
				12'd1700	: data2 <= weights[1701];
				12'd1701	: data2 <= weights[1702];
				12'd1702	: data2 <= weights[1703];
				12'd1703	: data2 <= weights[1704];
				12'd1704	: data2 <= weights[1705];
				12'd1705	: data2 <= weights[1706];
				12'd1706	: data2 <= weights[1707];
				12'd1707	: data2 <= weights[1708];
				12'd1708	: data2 <= weights[1709];
				12'd1709	: data2 <= weights[1710];
				12'd1710	: data2 <= weights[1711];
				12'd1711	: data2 <= weights[1712];
				12'd1712	: data2 <= weights[1713];
				12'd1713	: data2 <= weights[1714];
				12'd1714	: data2 <= weights[1715];
				12'd1715	: data2 <= weights[1716];
				12'd1716	: data2 <= weights[1717];
				12'd1717	: data2 <= weights[1718];
				12'd1718	: data2 <= weights[1719];
				12'd1719	: data2 <= weights[1720];
				12'd1720	: data2 <= weights[1721];
				12'd1721	: data2 <= weights[1722];
				12'd1722	: data2 <= weights[1723];
				12'd1723	: data2 <= weights[1724];
				12'd1724	: data2 <= weights[1725];
				12'd1725	: data2 <= weights[1726];
				12'd1726	: data2 <= weights[1727];
				12'd1727	: data2 <= weights[1728];
				12'd1728	: data2 <= weights[1729];
				12'd1729	: data2 <= weights[1730];
				12'd1730	: data2 <= weights[1731];
				12'd1731	: data2 <= weights[1732];
				12'd1732	: data2 <= weights[1733];
				12'd1733	: data2 <= weights[1734];
				12'd1734	: data2 <= weights[1735];
				12'd1735	: data2 <= weights[1736];
				12'd1736	: data2 <= weights[1737];
				12'd1737	: data2 <= weights[1738];
				12'd1738	: data2 <= weights[1739];
				12'd1739	: data2 <= weights[1740];
				12'd1740	: data2 <= weights[1741];
				12'd1741	: data2 <= weights[1742];
				12'd1742	: data2 <= weights[1743];
				12'd1743	: data2 <= weights[1744];
				12'd1744	: data2 <= weights[1745];
				12'd1745	: data2 <= weights[1746];
				12'd1746	: data2 <= weights[1747];
				12'd1747	: data2 <= weights[1748];
				12'd1748	: data2 <= weights[1749];
				12'd1749	: data2 <= weights[1750];
				12'd1750	: data2 <= weights[1751];
				12'd1751	: data2 <= weights[1752];
				12'd1752	: data2 <= weights[1753];
				12'd1753	: data2 <= weights[1754];
				12'd1754	: data2 <= weights[1755];
				12'd1755	: data2 <= weights[1756];
				12'd1756	: data2 <= weights[1757];
				12'd1757	: data2 <= weights[1758];
				12'd1758	: data2 <= weights[1759];
				12'd1759	: data2 <= weights[1760];
				12'd1760	: data2 <= weights[1761];
				12'd1761	: data2 <= weights[1762];
				12'd1762	: data2 <= weights[1763];
				12'd1763	: data2 <= weights[1764];
				12'd1764	: data2 <= weights[1765];
				12'd1765	: data2 <= weights[1766];
				12'd1766	: data2 <= weights[1767];
				12'd1767	: data2 <= weights[1768];
				12'd1768	: data2 <= weights[1769];
				12'd1769	: data2 <= weights[1770];
				12'd1770	: data2 <= weights[1771];
				12'd1771	: data2 <= weights[1772];
				12'd1772	: data2 <= weights[1773];
				12'd1773	: data2 <= weights[1774];
				12'd1774	: data2 <= weights[1775];
				12'd1775	: data2 <= weights[1776];
				12'd1776	: data2 <= weights[1777];
				12'd1777	: data2 <= weights[1778];
				12'd1778	: data2 <= weights[1779];
				12'd1779	: data2 <= weights[1780];
				12'd1780	: data2 <= weights[1781];
				12'd1781	: data2 <= weights[1782];
				12'd1782	: data2 <= weights[1783];
				12'd1783	: data2 <= weights[1784];
				12'd1784	: data2 <= weights[1785];
				12'd1785	: data2 <= weights[1786];
				12'd1786	: data2 <= weights[1787];
				12'd1787	: data2 <= weights[1788];
				12'd1788	: data2 <= weights[1789];
				12'd1789	: data2 <= weights[1790];
				12'd1790	: data2 <= weights[1791];
				12'd1791	: data2 <= weights[1792];
				12'd1792	: data2 <= weights[1793];
				12'd1793	: data2 <= weights[1794];
				12'd1794	: data2 <= weights[1795];
				12'd1795	: data2 <= weights[1796];
				12'd1796	: data2 <= weights[1797];
				12'd1797	: data2 <= weights[1798];
				12'd1798	: data2 <= weights[1799];
				12'd1799	: data2 <= weights[1800];
				12'd1800	: data2 <= weights[1801];
				12'd1801	: data2 <= weights[1802];
				12'd1802	: data2 <= weights[1803];
				12'd1803	: data2 <= weights[1804];
				12'd1804	: data2 <= weights[1805];
				12'd1805	: data2 <= weights[1806];
				12'd1806	: data2 <= weights[1807];
				12'd1807	: data2 <= weights[1808];
				12'd1808	: data2 <= weights[1809];
				12'd1809	: data2 <= weights[1810];
				12'd1810	: data2 <= weights[1811];
				12'd1811	: data2 <= weights[1812];
				12'd1812	: data2 <= weights[1813];
				12'd1813	: data2 <= weights[1814];
				12'd1814	: data2 <= weights[1815];
				12'd1815	: data2 <= weights[1816];
				12'd1816	: data2 <= weights[1817];
				12'd1817	: data2 <= weights[1818];
				12'd1818	: data2 <= weights[1819];
				12'd1819	: data2 <= weights[1820];
				12'd1820	: data2 <= weights[1821];
				12'd1821	: data2 <= weights[1822];
				12'd1822	: data2 <= weights[1823];
				12'd1823	: data2 <= weights[1824];
				12'd1824	: data2 <= weights[1825];
				12'd1825	: data2 <= weights[1826];
				12'd1826	: data2 <= weights[1827];
				12'd1827	: data2 <= weights[1828];
				12'd1828	: data2 <= weights[1829];
				12'd1829	: data2 <= weights[1830];
				12'd1830	: data2 <= weights[1831];
				12'd1831	: data2 <= weights[1832];
				12'd1832	: data2 <= weights[1833];
				12'd1833	: data2 <= weights[1834];
				12'd1834	: data2 <= weights[1835];
				12'd1835	: data2 <= weights[1836];
				12'd1836	: data2 <= weights[1837];
				12'd1837	: data2 <= weights[1838];
				12'd1838	: data2 <= weights[1839];
				12'd1839	: data2 <= weights[1840];
				12'd1840	: data2 <= weights[1841];
				12'd1841	: data2 <= weights[1842];
				12'd1842	: data2 <= weights[1843];
				12'd1843	: data2 <= weights[1844];
				12'd1844	: data2 <= weights[1845];
				12'd1845	: data2 <= weights[1846];
				12'd1846	: data2 <= weights[1847];
				12'd1847	: data2 <= weights[1848];
				12'd1848	: data2 <= weights[1849];
				12'd1849	: data2 <= weights[1850];
				12'd1850	: data2 <= weights[1851];
				12'd1851	: data2 <= weights[1852];
				12'd1852	: data2 <= weights[1853];
				12'd1853	: data2 <= weights[1854];
				12'd1854	: data2 <= weights[1855];
				12'd1855	: data2 <= weights[1856];
				12'd1856	: data2 <= weights[1857];
				12'd1857	: data2 <= weights[1858];
				12'd1858	: data2 <= weights[1859];
				12'd1859	: data2 <= weights[1860];
				12'd1860	: data2 <= weights[1861];
				12'd1861	: data2 <= weights[1862];
				12'd1862	: data2 <= weights[1863];
				12'd1863	: data2 <= weights[1864];
				12'd1864	: data2 <= weights[1865];
				12'd1865	: data2 <= weights[1866];
				12'd1866	: data2 <= weights[1867];
				12'd1867	: data2 <= weights[1868];
				12'd1868	: data2 <= weights[1869];
				12'd1869	: data2 <= weights[1870];
				12'd1870	: data2 <= weights[1871];
				12'd1871	: data2 <= weights[1872];
				12'd1872	: data2 <= weights[1873];
				12'd1873	: data2 <= weights[1874];
				12'd1874	: data2 <= weights[1875];
				12'd1875	: data2 <= weights[1876];
				12'd1876	: data2 <= weights[1877];
				12'd1877	: data2 <= weights[1878];
				12'd1878	: data2 <= weights[1879];
				12'd1879	: data2 <= weights[1880];
				12'd1880	: data2 <= weights[1881];
				12'd1881	: data2 <= weights[1882];
				12'd1882	: data2 <= weights[1883];
				12'd1883	: data2 <= weights[1884];
				12'd1884	: data2 <= weights[1885];
				12'd1885	: data2 <= weights[1886];
				12'd1886	: data2 <= weights[1887];
				12'd1887	: data2 <= weights[1888];
				12'd1888	: data2 <= weights[1889];
				12'd1889	: data2 <= weights[1890];
				12'd1890	: data2 <= weights[1891];
				12'd1891	: data2 <= weights[1892];
				12'd1892	: data2 <= weights[1893];
				12'd1893	: data2 <= weights[1894];
				12'd1894	: data2 <= weights[1895];
				12'd1895	: data2 <= weights[1896];
				12'd1896	: data2 <= weights[1897];
				12'd1897	: data2 <= weights[1898];
				12'd1898	: data2 <= weights[1899];
				12'd1899	: data2 <= weights[1900];
				12'd1900	: data2 <= weights[1901];
				12'd1901	: data2 <= weights[1902];
				12'd1902	: data2 <= weights[1903];
				12'd1903	: data2 <= weights[1904];
				12'd1904	: data2 <= weights[1905];
				12'd1905	: data2 <= weights[1906];
				12'd1906	: data2 <= weights[1907];
				12'd1907	: data2 <= weights[1908];
				12'd1908	: data2 <= weights[1909];
				12'd1909	: data2 <= weights[1910];
				12'd1910	: data2 <= weights[1911];
				12'd1911	: data2 <= weights[1912];
				12'd1912	: data2 <= weights[1913];
				12'd1913	: data2 <= weights[1914];
				12'd1914	: data2 <= weights[1915];
				12'd1915	: data2 <= weights[1916];
				12'd1916	: data2 <= weights[1917];
				12'd1917	: data2 <= weights[1918];
				12'd1918	: data2 <= weights[1919];
				12'd1919	: data2 <= weights[1920];
				12'd1920	: data2 <= weights[1921];
				12'd1921	: data2 <= weights[1922];
				12'd1922	: data2 <= weights[1923];
				12'd1923	: data2 <= weights[1924];
				12'd1924	: data2 <= weights[1925];
				12'd1925	: data2 <= weights[1926];
				12'd1926	: data2 <= weights[1927];
				12'd1927	: data2 <= weights[1928];
				12'd1928	: data2 <= weights[1929];
				12'd1929	: data2 <= weights[1930];
				12'd1930	: data2 <= weights[1931];
				12'd1931	: data2 <= weights[1932];
				12'd1932	: data2 <= weights[1933];
				12'd1933	: data2 <= weights[1934];
				12'd1934	: data2 <= weights[1935];
				12'd1935	: data2 <= weights[1936];
				12'd1936	: data2 <= weights[1937];
				12'd1937	: data2 <= weights[1938];
				12'd1938	: data2 <= weights[1939];
				12'd1939	: data2 <= weights[1940];
				12'd1940	: data2 <= weights[1941];
				12'd1941	: data2 <= weights[1942];
				12'd1942	: data2 <= weights[1943];
				12'd1943	: data2 <= weights[1944];
				12'd1944	: data2 <= weights[1945];
				12'd1945	: data2 <= weights[1946];
				12'd1946	: data2 <= weights[1947];
				12'd1947	: data2 <= weights[1948];
				12'd1948	: data2 <= weights[1949];
				12'd1949	: data2 <= weights[1950];
				12'd1950	: data2 <= weights[1951];
				12'd1951	: data2 <= weights[1952];
				12'd1952	: data2 <= weights[1953];
				12'd1953	: data2 <= weights[1954];
				12'd1954	: data2 <= weights[1955];
				12'd1955	: data2 <= weights[1956];
				12'd1956	: data2 <= weights[1957];
				12'd1957	: data2 <= weights[1958];
				12'd1958	: data2 <= weights[1959];
				12'd1959	: data2 <= weights[1960];
				12'd1960	: data2 <= weights[1961];
				12'd1961	: data2 <= weights[1962];
				12'd1962	: data2 <= weights[1963];
				12'd1963	: data2 <= weights[1964];
				12'd1964	: data2 <= weights[1965];
				12'd1965	: data2 <= weights[1966];
				12'd1966	: data2 <= weights[1967];
				12'd1967	: data2 <= weights[1968];
				12'd1968	: data2 <= weights[1969];
				12'd1969	: data2 <= weights[1970];
				12'd1970	: data2 <= weights[1971];
				12'd1971	: data2 <= weights[1972];
				12'd1972	: data2 <= weights[1973];
				12'd1973	: data2 <= weights[1974];
				12'd1974	: data2 <= weights[1975];
				12'd1975	: data2 <= weights[1976];
				12'd1976	: data2 <= weights[1977];
				12'd1977	: data2 <= weights[1978];
				12'd1978	: data2 <= weights[1979];
				12'd1979	: data2 <= weights[1980];
				12'd1980	: data2 <= weights[1981];
				12'd1981	: data2 <= weights[1982];
				12'd1982	: data2 <= weights[1983];
				12'd1983	: data2 <= weights[1984];
				12'd1984	: data2 <= weights[1985];
				12'd1985	: data2 <= weights[1986];
				12'd1986	: data2 <= weights[1987];
				12'd1987	: data2 <= weights[1988];
				12'd1988	: data2 <= weights[1989];
				12'd1989	: data2 <= weights[1990];
				12'd1990	: data2 <= weights[1991];
				12'd1991	: data2 <= weights[1992];
				12'd1992	: data2 <= weights[1993];
				12'd1993	: data2 <= weights[1994];
				12'd1994	: data2 <= weights[1995];
				12'd1995	: data2 <= weights[1996];
				12'd1996	: data2 <= weights[1997];
				12'd1997	: data2 <= weights[1998];
				12'd1998	: data2 <= weights[1999];
				12'd1999	: data2 <= weights[2000];
				12'd2000	: data2 <= weights[2001];
				12'd2001	: data2 <= weights[2002];
				12'd2002	: data2 <= weights[2003];
				12'd2003	: data2 <= weights[2004];
				12'd2004	: data2 <= weights[2005];
				12'd2005	: data2 <= weights[2006];
				12'd2006	: data2 <= weights[2007];
				12'd2007	: data2 <= weights[2008];
				12'd2008	: data2 <= weights[2009];
				12'd2009	: data2 <= weights[2010];
				12'd2010	: data2 <= weights[2011];
				12'd2011	: data2 <= weights[2012];
				12'd2012	: data2 <= weights[2013];
				12'd2013	: data2 <= weights[2014];
				12'd2014	: data2 <= weights[2015];
				12'd2015	: data2 <= weights[2016];
				12'd2016	: data2 <= weights[2017];
				12'd2017	: data2 <= weights[2018];
				12'd2018	: data2 <= weights[2019];
				12'd2019	: data2 <= weights[2020];
				12'd2020	: data2 <= weights[2021];
				12'd2021	: data2 <= weights[2022];
				12'd2022	: data2 <= weights[2023];
				12'd2023	: data2 <= weights[2024];
				12'd2024	: data2 <= weights[2025];
				12'd2025	: data2 <= weights[2026];
				12'd2026	: data2 <= weights[2027];
				12'd2027	: data2 <= weights[2028];
				12'd2028	: data2 <= weights[2029];
				12'd2029	: data2 <= weights[2030];
				12'd2030	: data2 <= weights[2031];
				12'd2031	: data2 <= weights[2032];
				12'd2032	: data2 <= weights[2033];
				12'd2033	: data2 <= weights[2034];
				12'd2034	: data2 <= weights[2035];
				12'd2035	: data2 <= weights[2036];
				12'd2036	: data2 <= weights[2037];
				12'd2037	: data2 <= weights[2038];
				12'd2038	: data2 <= weights[2039];
				12'd2039	: data2 <= weights[2040];
				12'd2040	: data2 <= weights[2041];
				12'd2041	: data2 <= weights[2042];
				12'd2042	: data2 <= weights[2043];
				12'd2043	: data2 <= weights[2044];
				12'd2044	: data2 <= weights[2045];
				12'd2045	: data2 <= weights[2046];
				12'd2046	: data2 <= weights[2047];
				12'd2047	: data2 <= weights[2048];
				12'd2048	: data2 <= weights[2049];
				12'd2049	: data2 <= weights[2050];
				12'd2050	: data2 <= weights[2051];
				12'd2051	: data2 <= weights[2052];
				12'd2052	: data2 <= weights[2053];
				12'd2053	: data2 <= weights[2054];
				12'd2054	: data2 <= weights[2055];
				12'd2055	: data2 <= weights[2056];
				12'd2056	: data2 <= weights[2057];
				12'd2057	: data2 <= weights[2058];
				12'd2058	: data2 <= weights[2059];
				12'd2059	: data2 <= weights[2060];
				12'd2060	: data2 <= weights[2061];
				12'd2061	: data2 <= weights[2062];
				12'd2062	: data2 <= weights[2063];
				12'd2063	: data2 <= weights[2064];
				12'd2064	: data2 <= weights[2065];
				12'd2065	: data2 <= weights[2066];
				12'd2066	: data2 <= weights[2067];
				12'd2067	: data2 <= weights[2068];
				12'd2068	: data2 <= weights[2069];
				12'd2069	: data2 <= weights[2070];
				12'd2070	: data2 <= weights[2071];
				12'd2071	: data2 <= weights[2072];
				12'd2072	: data2 <= weights[2073];
				12'd2073	: data2 <= weights[2074];
				12'd2074	: data2 <= weights[2075];
				12'd2075	: data2 <= weights[2076];
				12'd2076	: data2 <= weights[2077];
				12'd2077	: data2 <= weights[2078];
				12'd2078	: data2 <= weights[2079];
				12'd2079	: data2 <= weights[2080];
				12'd2080	: data2 <= weights[2081];
				12'd2081	: data2 <= weights[2082];
				12'd2082	: data2 <= weights[2083];
				12'd2083	: data2 <= weights[2084];
				12'd2084	: data2 <= weights[2085];
				12'd2085	: data2 <= weights[2086];
				12'd2086	: data2 <= weights[2087];
				12'd2087	: data2 <= weights[2088];
				12'd2088	: data2 <= weights[2089];
				12'd2089	: data2 <= weights[2090];
				12'd2090	: data2 <= weights[2091];
				12'd2091	: data2 <= weights[2092];
				12'd2092	: data2 <= weights[2093];
				12'd2093	: data2 <= weights[2094];
				12'd2094	: data2 <= weights[2095];
				12'd2095	: data2 <= weights[2096];
				12'd2096	: data2 <= weights[2097];
				12'd2097	: data2 <= weights[2098];
				12'd2098	: data2 <= weights[2099];
				12'd2099	: data2 <= weights[2100];
				12'd2100	: data2 <= weights[2101];
				12'd2101	: data2 <= weights[2102];
				12'd2102	: data2 <= weights[2103];
				12'd2103	: data2 <= weights[2104];
				12'd2104	: data2 <= weights[2105];
				12'd2105	: data2 <= weights[2106];
				12'd2106	: data2 <= weights[2107];
				12'd2107	: data2 <= weights[2108];
				12'd2108	: data2 <= weights[2109];
				12'd2109	: data2 <= weights[2110];
				12'd2110	: data2 <= weights[2111];
				12'd2111	: data2 <= weights[2112];
				12'd2112	: data2 <= weights[2113];
				12'd2113	: data2 <= weights[2114];
				12'd2114	: data2 <= weights[2115];
				12'd2115	: data2 <= weights[2116];
				12'd2116	: data2 <= weights[2117];
				12'd2117	: data2 <= weights[2118];
				12'd2118	: data2 <= weights[2119];
				12'd2119	: data2 <= weights[2120];
				12'd2120	: data2 <= weights[2121];
				12'd2121	: data2 <= weights[2122];
				12'd2122	: data2 <= weights[2123];
				12'd2123	: data2 <= weights[2124];
				12'd2124	: data2 <= weights[2125];
				12'd2125	: data2 <= weights[2126];
				12'd2126	: data2 <= weights[2127];
				12'd2127	: data2 <= weights[2128];
				12'd2128	: data2 <= weights[2129];
				12'd2129	: data2 <= weights[2130];
				12'd2130	: data2 <= weights[2131];
				12'd2131	: data2 <= weights[2132];
				12'd2132	: data2 <= weights[2133];
				12'd2133	: data2 <= weights[2134];
				12'd2134	: data2 <= weights[2135];
				12'd2135	: data2 <= weights[2136];
				12'd2136	: data2 <= weights[2137];
				12'd2137	: data2 <= weights[2138];
				12'd2138	: data2 <= weights[2139];
				12'd2139	: data2 <= weights[2140];
				12'd2140	: data2 <= weights[2141];
				12'd2141	: data2 <= weights[2142];
				12'd2142	: data2 <= weights[2143];
				12'd2143	: data2 <= weights[2144];
				12'd2144	: data2 <= weights[2145];
				12'd2145	: data2 <= weights[2146];
				12'd2146	: data2 <= weights[2147];
				12'd2147	: data2 <= weights[2148];
				12'd2148	: data2 <= weights[2149];
				12'd2149	: data2 <= weights[2150];
				12'd2150	: data2 <= weights[2151];
				12'd2151	: data2 <= weights[2152];
				12'd2152	: data2 <= weights[2153];
				12'd2153	: data2 <= weights[2154];
				12'd2154	: data2 <= weights[2155];
				12'd2155	: data2 <= weights[2156];
				12'd2156	: data2 <= weights[2157];
				12'd2157	: data2 <= weights[2158];
				12'd2158	: data2 <= weights[2159];
				12'd2159	: data2 <= weights[2160];
				12'd2160	: data2 <= weights[2161];
				12'd2161	: data2 <= weights[2162];
				12'd2162	: data2 <= weights[2163];
				12'd2163	: data2 <= weights[2164];
				12'd2164	: data2 <= weights[2165];
				12'd2165	: data2 <= weights[2166];
				12'd2166	: data2 <= weights[2167];
				12'd2167	: data2 <= weights[2168];
				12'd2168	: data2 <= weights[2169];
				12'd2169	: data2 <= weights[2170];
				12'd2170	: data2 <= weights[2171];
				12'd2171	: data2 <= weights[2172];
				12'd2172	: data2 <= weights[2173];
				12'd2173	: data2 <= weights[2174];
				12'd2174	: data2 <= weights[2175];
				12'd2175	: data2 <= weights[2176];
				12'd2176	: data2 <= weights[2177];
				12'd2177	: data2 <= weights[2178];
				12'd2178	: data2 <= weights[2179];
				12'd2179	: data2 <= weights[2180];
				12'd2180	: data2 <= weights[2181];
				12'd2181	: data2 <= weights[2182];
				12'd2182	: data2 <= weights[2183];
				12'd2183	: data2 <= weights[2184];
				12'd2184	: data2 <= weights[2185];
				12'd2185	: data2 <= weights[2186];
				12'd2186	: data2 <= weights[2187];
				12'd2187	: data2 <= weights[2188];
				12'd2188	: data2 <= weights[2189];
				12'd2189	: data2 <= weights[2190];
				12'd2190	: data2 <= weights[2191];
				12'd2191	: data2 <= weights[2192];
				12'd2192	: data2 <= weights[2193];
				12'd2193	: data2 <= weights[2194];
				12'd2194	: data2 <= weights[2195];
				12'd2195	: data2 <= weights[2196];
				12'd2196	: data2 <= weights[2197];
				12'd2197	: data2 <= weights[2198];
				12'd2198	: data2 <= weights[2199];
				12'd2199	: data2 <= weights[2200];
				12'd2200	: data2 <= weights[2201];
				12'd2201	: data2 <= weights[2202];
				12'd2202	: data2 <= weights[2203];
				12'd2203	: data2 <= weights[2204];
				12'd2204	: data2 <= weights[2205];
				12'd2205	: data2 <= weights[2206];
				12'd2206	: data2 <= weights[2207];
				12'd2207	: data2 <= weights[2208];
				12'd2208	: data2 <= weights[2209];
				12'd2209	: data2 <= weights[2210];
				12'd2210	: data2 <= weights[2211];
				12'd2211	: data2 <= weights[2212];
				12'd2212	: data2 <= weights[2213];
				12'd2213	: data2 <= weights[2214];
				12'd2214	: data2 <= weights[2215];
				12'd2215	: data2 <= weights[2216];
				12'd2216	: data2 <= weights[2217];
				12'd2217	: data2 <= weights[2218];
				12'd2218	: data2 <= weights[2219];
				12'd2219	: data2 <= weights[2220];
				12'd2220	: data2 <= weights[2221];
				12'd2221	: data2 <= weights[2222];
				12'd2222	: data2 <= weights[2223];
				12'd2223	: data2 <= weights[2224];
				12'd2224	: data2 <= weights[2225];
				12'd2225	: data2 <= weights[2226];
				12'd2226	: data2 <= weights[2227];
				12'd2227	: data2 <= weights[2228];
				12'd2228	: data2 <= weights[2229];
				12'd2229	: data2 <= weights[2230];
				12'd2230	: data2 <= weights[2231];
				12'd2231	: data2 <= weights[2232];
				12'd2232	: data2 <= weights[2233];
				12'd2233	: data2 <= weights[2234];
				12'd2234	: data2 <= weights[2235];
				12'd2235	: data2 <= weights[2236];
				12'd2236	: data2 <= weights[2237];
				12'd2237	: data2 <= weights[2238];
				12'd2238	: data2 <= weights[2239];
				12'd2239	: data2 <= weights[2240];
				12'd2240	: data2 <= weights[2241];
				12'd2241	: data2 <= weights[2242];
				12'd2242	: data2 <= weights[2243];
				12'd2243	: data2 <= weights[2244];
				12'd2244	: data2 <= weights[2245];
				12'd2245	: data2 <= weights[2246];
				12'd2246	: data2 <= weights[2247];
				12'd2247	: data2 <= weights[2248];
				12'd2248	: data2 <= weights[2249];
				12'd2249	: data2 <= weights[2250];
				12'd2250	: data2 <= weights[2251];
				12'd2251	: data2 <= weights[2252];
				12'd2252	: data2 <= weights[2253];
				12'd2253	: data2 <= weights[2254];
				12'd2254	: data2 <= weights[2255];
				12'd2255	: data2 <= weights[2256];
				12'd2256	: data2 <= weights[2257];
				12'd2257	: data2 <= weights[2258];
				12'd2258	: data2 <= weights[2259];
				12'd2259	: data2 <= weights[2260];
				12'd2260	: data2 <= weights[2261];
				12'd2261	: data2 <= weights[2262];
				12'd2262	: data2 <= weights[2263];
				12'd2263	: data2 <= weights[2264];
				12'd2264	: data2 <= weights[2265];
				12'd2265	: data2 <= weights[2266];
				12'd2266	: data2 <= weights[2267];
				12'd2267	: data2 <= weights[2268];
				12'd2268	: data2 <= weights[2269];
				12'd2269	: data2 <= weights[2270];
				12'd2270	: data2 <= weights[2271];
				12'd2271	: data2 <= weights[2272];
				12'd2272	: data2 <= weights[2273];
				12'd2273	: data2 <= weights[2274];
				12'd2274	: data2 <= weights[2275];
				12'd2275	: data2 <= weights[2276];
				12'd2276	: data2 <= weights[2277];
				12'd2277	: data2 <= weights[2278];
				12'd2278	: data2 <= weights[2279];
				12'd2279	: data2 <= weights[2280];
				12'd2280	: data2 <= weights[2281];
				12'd2281	: data2 <= weights[2282];
				12'd2282	: data2 <= weights[2283];
				12'd2283	: data2 <= weights[2284];
				12'd2284	: data2 <= weights[2285];
				12'd2285	: data2 <= weights[2286];
				12'd2286	: data2 <= weights[2287];
				12'd2287	: data2 <= weights[2288];
				12'd2288	: data2 <= weights[2289];
				12'd2289	: data2 <= weights[2290];
				12'd2290	: data2 <= weights[2291];
				12'd2291	: data2 <= weights[2292];
				12'd2292	: data2 <= weights[2293];
				12'd2293	: data2 <= weights[2294];
				12'd2294	: data2 <= weights[2295];
				12'd2295	: data2 <= weights[2296];
				12'd2296	: data2 <= weights[2297];
				12'd2297	: data2 <= weights[2298];
				12'd2298	: data2 <= weights[2299];
				12'd2299	: data2 <= weights[2300];
				12'd2300	: data2 <= weights[2301];
				12'd2301	: data2 <= weights[2302];
				12'd2302	: data2 <= weights[2303];
				12'd2303	: data2 <= weights[2304];
				12'd2304	: data2 <= weights[2305];
				12'd2305	: data2 <= weights[2306];
				12'd2306	: data2 <= weights[2307];
				12'd2307	: data2 <= weights[2308];
				12'd2308	: data2 <= weights[2309];
				12'd2309	: data2 <= weights[2310];
				12'd2310	: data2 <= weights[2311];
				12'd2311	: data2 <= weights[2312];
				12'd2312	: data2 <= weights[2313];
				12'd2313	: data2 <= weights[2314];
				12'd2314	: data2 <= weights[2315];
				12'd2315	: data2 <= weights[2316];
				12'd2316	: data2 <= weights[2317];
				12'd2317	: data2 <= weights[2318];
				12'd2318	: data2 <= weights[2319];
				12'd2319	: data2 <= weights[2320];
				12'd2320	: data2 <= weights[2321];
				12'd2321	: data2 <= weights[2322];
				12'd2322	: data2 <= weights[2323];
				12'd2323	: data2 <= weights[2324];
				12'd2324	: data2 <= weights[2325];
				12'd2325	: data2 <= weights[2326];
				12'd2326	: data2 <= weights[2327];
				12'd2327	: data2 <= weights[2328];
				12'd2328	: data2 <= weights[2329];
				12'd2329	: data2 <= weights[2330];
				12'd2330	: data2 <= weights[2331];
				12'd2331	: data2 <= weights[2332];
				12'd2332	: data2 <= weights[2333];
				12'd2333	: data2 <= weights[2334];
				12'd2334	: data2 <= weights[2335];
				12'd2335	: data2 <= weights[2336];
				12'd2336	: data2 <= weights[2337];
				12'd2337	: data2 <= weights[2338];
				12'd2338	: data2 <= weights[2339];
				12'd2339	: data2 <= weights[2340];
				12'd2340	: data2 <= weights[2341];
				12'd2341	: data2 <= weights[2342];
				12'd2342	: data2 <= weights[2343];
				12'd2343	: data2 <= weights[2344];
				12'd2344	: data2 <= weights[2345];
				12'd2345	: data2 <= weights[2346];
				12'd2346	: data2 <= weights[2347];
				12'd2347	: data2 <= weights[2348];
				12'd2348	: data2 <= weights[2349];
				12'd2349	: data2 <= weights[2350];
				12'd2350	: data2 <= weights[2351];
				12'd2351	: data2 <= weights[2352];
				12'd2352	: data2 <= weights[2353];
				12'd2353	: data2 <= weights[2354];
				12'd2354	: data2 <= weights[2355];
				12'd2355	: data2 <= weights[2356];
				12'd2356	: data2 <= weights[2357];
				12'd2357	: data2 <= weights[2358];
				12'd2358	: data2 <= weights[2359];
				12'd2359	: data2 <= weights[2360];
				12'd2360	: data2 <= weights[2361];
				12'd2361	: data2 <= weights[2362];
				12'd2362	: data2 <= weights[2363];
				12'd2363	: data2 <= weights[2364];
				12'd2364	: data2 <= weights[2365];
				12'd2365	: data2 <= weights[2366];
				12'd2366	: data2 <= weights[2367];
				12'd2367	: data2 <= weights[2368];
				12'd2368	: data2 <= weights[2369];
				12'd2369	: data2 <= weights[2370];
				12'd2370	: data2 <= weights[2371];
				12'd2371	: data2 <= weights[2372];
				12'd2372	: data2 <= weights[2373];
				12'd2373	: data2 <= weights[2374];
				12'd2374	: data2 <= weights[2375];
				12'd2375	: data2 <= weights[2376];
				12'd2376	: data2 <= weights[2377];
				12'd2377	: data2 <= weights[2378];
				12'd2378	: data2 <= weights[2379];
				12'd2379	: data2 <= weights[2380];
				12'd2380	: data2 <= weights[2381];
				12'd2381	: data2 <= weights[2382];
				12'd2382	: data2 <= weights[2383];
				12'd2383	: data2 <= weights[2384];
				12'd2384	: data2 <= weights[2385];
				12'd2385	: data2 <= weights[2386];
				12'd2386	: data2 <= weights[2387];
				12'd2387	: data2 <= weights[2388];
				12'd2388	: data2 <= weights[2389];
				12'd2389	: data2 <= weights[2390];
				12'd2390	: data2 <= weights[2391];
				12'd2391	: data2 <= weights[2392];
				12'd2392	: data2 <= weights[2393];
				12'd2393	: data2 <= weights[2394];
				12'd2394	: data2 <= weights[2395];
				12'd2395	: data2 <= weights[2396];
				12'd2396	: data2 <= weights[2397];
				12'd2397	: data2 <= weights[2398];
				12'd2398	: data2 <= weights[2399];
				12'd2399	: data2 <= weights[2400];
				12'd2400	: data2 <= weights[2401];
				12'd2401	: data2 <= weights[2402];
				12'd2402	: data2 <= weights[2403];
				12'd2403	: data2 <= weights[2404];
				12'd2404	: data2 <= weights[2405];
				12'd2405	: data2 <= weights[2406];
				12'd2406	: data2 <= weights[2407];
				12'd2407	: data2 <= weights[2408];
				12'd2408	: data2 <= weights[2409];
				12'd2409	: data2 <= weights[2410];
				12'd2410	: data2 <= weights[2411];
				12'd2411	: data2 <= weights[2412];
				12'd2412	: data2 <= weights[2413];
				12'd2413	: data2 <= weights[2414];
				12'd2414	: data2 <= weights[2415];
				12'd2415	: data2 <= weights[2416];
				12'd2416	: data2 <= weights[2417];
				12'd2417	: data2 <= weights[2418];
				12'd2418	: data2 <= weights[2419];
				12'd2419	: data2 <= weights[2420];
				12'd2420	: data2 <= weights[2421];
				12'd2421	: data2 <= weights[2422];
				12'd2422	: data2 <= weights[2423];
				12'd2423	: data2 <= weights[2424];
				12'd2424	: data2 <= weights[2425];
				12'd2425	: data2 <= weights[2426];
				12'd2426	: data2 <= weights[2427];
				12'd2427	: data2 <= weights[2428];
				12'd2428	: data2 <= weights[2429];
				12'd2429	: data2 <= weights[2430];
				12'd2430	: data2 <= weights[2431];
				12'd2431	: data2 <= weights[2432];
				12'd2432	: data2 <= weights[2433];
				12'd2433	: data2 <= weights[2434];
				12'd2434	: data2 <= weights[2435];
				12'd2435	: data2 <= weights[2436];
				12'd2436	: data2 <= weights[2437];
				12'd2437	: data2 <= weights[2438];
				12'd2438	: data2 <= weights[2439];
				12'd2439	: data2 <= weights[2440];
				12'd2440	: data2 <= weights[2441];
				12'd2441	: data2 <= weights[2442];
				12'd2442	: data2 <= weights[2443];
				12'd2443	: data2 <= weights[2444];
				12'd2444	: data2 <= weights[2445];
				12'd2445	: data2 <= weights[2446];
				12'd2446	: data2 <= weights[2447];
				12'd2447	: data2 <= weights[2448];
				12'd2448	: data2 <= weights[2449];
				12'd2449	: data2 <= weights[2450];
				12'd2450	: data2 <= weights[2451];
				12'd2451	: data2 <= weights[2452];
				12'd2452	: data2 <= weights[2453];
				12'd2453	: data2 <= weights[2454];
				12'd2454	: data2 <= weights[2455];
				12'd2455	: data2 <= weights[2456];
				12'd2456	: data2 <= weights[2457];
				12'd2457	: data2 <= weights[2458];
				12'd2458	: data2 <= weights[2459];
				12'd2459	: data2 <= weights[2460];
				12'd2460	: data2 <= weights[2461];
				12'd2461	: data2 <= weights[2462];
				12'd2462	: data2 <= weights[2463];
				12'd2463	: data2 <= weights[2464];
				12'd2464	: data2 <= weights[2465];
				12'd2465	: data2 <= weights[2466];
				12'd2466	: data2 <= weights[2467];
				12'd2467	: data2 <= weights[2468];
				12'd2468	: data2 <= weights[2469];
				12'd2469	: data2 <= weights[2470];
				12'd2470	: data2 <= weights[2471];
				12'd2471	: data2 <= weights[2472];
				12'd2472	: data2 <= weights[2473];
				12'd2473	: data2 <= weights[2474];
				12'd2474	: data2 <= weights[2475];
				12'd2475	: data2 <= weights[2476];
				12'd2476	: data2 <= weights[2477];
				12'd2477	: data2 <= weights[2478];
				12'd2478	: data2 <= weights[2479];
				12'd2479	: data2 <= weights[2480];
				12'd2480	: data2 <= weights[2481];
				12'd2481	: data2 <= weights[2482];
				12'd2482	: data2 <= weights[2483];
				12'd2483	: data2 <= weights[2484];
				12'd2484	: data2 <= weights[2485];
				12'd2485	: data2 <= weights[2486];
				12'd2486	: data2 <= weights[2487];
				12'd2487	: data2 <= weights[2488];
				12'd2488	: data2 <= weights[2489];
				12'd2489	: data2 <= weights[2490];
				12'd2490	: data2 <= weights[2491];
				12'd2491	: data2 <= weights[2492];
				12'd2492	: data2 <= weights[2493];
				12'd2493	: data2 <= weights[2494];
				12'd2494	: data2 <= weights[2495];
				12'd2495	: data2 <= weights[2496];
				12'd2496	: data2 <= weights[2497];
				12'd2497	: data2 <= weights[2498];
				12'd2498	: data2 <= weights[2499];
				12'd2499	: data2 <= weights[2500];
				12'd2500	: data2 <= weights[2501];
				12'd2501	: data2 <= weights[2502];
				12'd2502	: data2 <= weights[2503];
				12'd2503	: data2 <= weights[2504];
				12'd2504	: data2 <= weights[2505];
				12'd2505	: data2 <= weights[2506];
				12'd2506	: data2 <= weights[2507];
				12'd2507	: data2 <= weights[2508];
				12'd2508	: data2 <= weights[2509];
				12'd2509	: data2 <= weights[2510];
				12'd2510	: data2 <= weights[2511];
				12'd2511	: data2 <= weights[2512];
				12'd2512	: data2 <= weights[2513];
				12'd2513	: data2 <= weights[2514];
				12'd2514	: data2 <= weights[2515];
				12'd2515	: data2 <= weights[2516];
				12'd2516	: data2 <= weights[2517];
				12'd2517	: data2 <= weights[2518];
				12'd2518	: data2 <= weights[2519];
				12'd2519	: data2 <= weights[2520];
				12'd2520	: data2 <= weights[2521];
				12'd2521	: data2 <= weights[2522];
				12'd2522	: data2 <= weights[2523];
				12'd2523	: data2 <= weights[2524];
				12'd2524	: data2 <= weights[2525];
				12'd2525	: data2 <= weights[2526];
				12'd2526	: data2 <= weights[2527];
				12'd2527	: data2 <= weights[2528];
				12'd2528	: data2 <= weights[2529];
				12'd2529	: data2 <= weights[2530];
				12'd2530	: data2 <= weights[2531];
				12'd2531	: data2 <= weights[2532];
				12'd2532	: data2 <= weights[2533];
				12'd2533	: data2 <= weights[2534];
				12'd2534	: data2 <= weights[2535];
				12'd2535	: data2 <= weights[2536];
				12'd2536	: data2 <= weights[2537];
				12'd2537	: data2 <= weights[2538];
				12'd2538	: data2 <= weights[2539];
				12'd2539	: data2 <= weights[2540];
				12'd2540	: data2 <= weights[2541];
				12'd2541	: data2 <= weights[2542];
				12'd2542	: data2 <= weights[2543];
				12'd2543	: data2 <= weights[2544];
				12'd2544	: data2 <= weights[2545];
				12'd2545	: data2 <= weights[2546];
				12'd2546	: data2 <= weights[2547];
				12'd2547	: data2 <= weights[2548];
				12'd2548	: data2 <= weights[2549];
				12'd2549	: data2 <= weights[2550];
				12'd2550	: data2 <= weights[2551];
				12'd2551	: data2 <= weights[2552];
				12'd2552	: data2 <= weights[2553];
				12'd2553	: data2 <= weights[2554];
				12'd2554	: data2 <= weights[2555];
				12'd2555	: data2 <= weights[2556];
				12'd2556	: data2 <= weights[2557];
				12'd2557	: data2 <= weights[2558];
				12'd2558	: data2 <= weights[2559];
				12'd2559	: data2 <= weights[2560];
				12'd2560	: data2 <= weights[2561];
				12'd2561	: data2 <= weights[2562];
				12'd2562	: data2 <= weights[2563];
				12'd2563	: data2 <= weights[2564];
				12'd2564	: data2 <= weights[2565];
				12'd2565	: data2 <= weights[2566];
				12'd2566	: data2 <= weights[2567];
				12'd2567	: data2 <= weights[2568];
				12'd2568	: data2 <= weights[2569];
				12'd2569	: data2 <= weights[2570];
				12'd2570	: data2 <= weights[2571];
				12'd2571	: data2 <= weights[2572];
				12'd2572	: data2 <= weights[2573];
				12'd2573	: data2 <= weights[2574];
				12'd2574	: data2 <= weights[2575];
				12'd2575	: data2 <= weights[2576];
				12'd2576	: data2 <= weights[2577];
				12'd2577	: data2 <= weights[2578];
				12'd2578	: data2 <= weights[2579];
				12'd2579	: data2 <= weights[2580];
				12'd2580	: data2 <= weights[2581];
				12'd2581	: data2 <= weights[2582];
				12'd2582	: data2 <= weights[2583];
				12'd2583	: data2 <= weights[2584];
				12'd2584	: data2 <= weights[2585];
				12'd2585	: data2 <= weights[2586];
				12'd2586	: data2 <= weights[2587];
				12'd2587	: data2 <= weights[2588];
				12'd2588	: data2 <= weights[2589];
				12'd2589	: data2 <= weights[2590];
				12'd2590	: data2 <= weights[2591];
				12'd2591	: data2 <= weights[2592];
				12'd2592	: data2 <= weights[2593];
				12'd2593	: data2 <= weights[2594];
				12'd2594	: data2 <= weights[2595];
				12'd2595	: data2 <= weights[2596];
				12'd2596	: data2 <= weights[2597];
				12'd2597	: data2 <= weights[2598];
				12'd2598	: data2 <= weights[2599];
				12'd2599	: data2 <= weights[2600];
				12'd2600	: data2 <= weights[2601];
				12'd2601	: data2 <= weights[2602];
				12'd2602	: data2 <= weights[2603];
				12'd2603	: data2 <= weights[2604];
				12'd2604	: data2 <= weights[2605];
				12'd2605	: data2 <= weights[2606];
				12'd2606	: data2 <= weights[2607];
				12'd2607	: data2 <= weights[2608];
				12'd2608	: data2 <= weights[2609];
				12'd2609	: data2 <= weights[2610];
				12'd2610	: data2 <= weights[2611];
				12'd2611	: data2 <= weights[2612];
				12'd2612	: data2 <= weights[2613];
				12'd2613	: data2 <= weights[2614];
				12'd2614	: data2 <= weights[2615];
				12'd2615	: data2 <= weights[2616];
				12'd2616	: data2 <= weights[2617];
				12'd2617	: data2 <= weights[2618];
				12'd2618	: data2 <= weights[2619];
				12'd2619	: data2 <= weights[2620];
				12'd2620	: data2 <= weights[2621];
				12'd2621	: data2 <= weights[2622];
				12'd2622	: data2 <= weights[2623];
				12'd2623	: data2 <= weights[2624];
				12'd2624	: data2 <= weights[2625];
				12'd2625	: data2 <= weights[2626];
				12'd2626	: data2 <= weights[2627];
				12'd2627	: data2 <= weights[2628];
				12'd2628	: data2 <= weights[2629];
				12'd2629	: data2 <= weights[2630];
				12'd2630	: data2 <= weights[2631];
				12'd2631	: data2 <= weights[2632];
				12'd2632	: data2 <= weights[2633];
				12'd2633	: data2 <= weights[2634];
				12'd2634	: data2 <= weights[2635];
				12'd2635	: data2 <= weights[2636];
				12'd2636	: data2 <= weights[2637];
				12'd2637	: data2 <= weights[2638];
				12'd2638	: data2 <= weights[2639];
				12'd2639	: data2 <= weights[2640];
				12'd2640	: data2 <= weights[2641];
				12'd2641	: data2 <= weights[2642];
				12'd2642	: data2 <= weights[2643];
				12'd2643	: data2 <= weights[2644];
				12'd2644	: data2 <= weights[2645];
				12'd2645	: data2 <= weights[2646];
				12'd2646	: data2 <= weights[2647];
				12'd2647	: data2 <= weights[2648];
				12'd2648	: data2 <= weights[2649];
				12'd2649	: data2 <= weights[2650];
				12'd2650	: data2 <= weights[2651];
				12'd2651	: data2 <= weights[2652];
				12'd2652	: data2 <= weights[2653];
				12'd2653	: data2 <= weights[2654];
				12'd2654	: data2 <= weights[2655];
				12'd2655	: data2 <= weights[2656];
				12'd2656	: data2 <= weights[2657];
				12'd2657	: data2 <= weights[2658];
				12'd2658	: data2 <= weights[2659];
				12'd2659	: data2 <= weights[2660];
				12'd2660	: data2 <= weights[2661];
				12'd2661	: data2 <= weights[2662];
				12'd2662	: data2 <= weights[2663];
				12'd2663	: data2 <= weights[2664];
				12'd2664	: data2 <= weights[2665];
				12'd2665	: data2 <= weights[2666];
				12'd2666	: data2 <= weights[2667];
				12'd2667	: data2 <= weights[2668];
				12'd2668	: data2 <= weights[2669];
				12'd2669	: data2 <= weights[2670];
				12'd2670	: data2 <= weights[2671];
				12'd2671	: data2 <= weights[2672];
				12'd2672	: data2 <= weights[2673];
				12'd2673	: data2 <= weights[2674];
				12'd2674	: data2 <= weights[2675];
				12'd2675	: data2 <= weights[2676];
				12'd2676	: data2 <= weights[2677];
				12'd2677	: data2 <= weights[2678];
				12'd2678	: data2 <= weights[2679];
				12'd2679	: data2 <= weights[2680];
				12'd2680	: data2 <= weights[2681];
				12'd2681	: data2 <= weights[2682];
				12'd2682	: data2 <= weights[2683];
				12'd2683	: data2 <= weights[2684];
				12'd2684	: data2 <= weights[2685];
				12'd2685	: data2 <= weights[2686];
				12'd2686	: data2 <= weights[2687];
				12'd2687	: data2 <= weights[2688];
				12'd2688	: data2 <= weights[2689];
				12'd2689	: data2 <= weights[2690];
				12'd2690	: data2 <= weights[2691];
				12'd2691	: data2 <= weights[2692];
				12'd2692	: data2 <= weights[2693];
				12'd2693	: data2 <= weights[2694];
				12'd2694	: data2 <= weights[2695];
				12'd2695	: data2 <= weights[2696];
				12'd2696	: data2 <= weights[2697];
				12'd2697	: data2 <= weights[2698];
				12'd2698	: data2 <= weights[2699];
				12'd2699	: data2 <= weights[2700];
				12'd2700	: data2 <= weights[2701];
				12'd2701	: data2 <= weights[2702];
				12'd2702	: data2 <= weights[2703];
				12'd2703	: data2 <= weights[2704];
				12'd2704	: data2 <= weights[2705];
				12'd2705	: data2 <= weights[2706];
				12'd2706	: data2 <= weights[2707];
				12'd2707	: data2 <= weights[2708];
				12'd2708	: data2 <= weights[2709];
				12'd2709	: data2 <= weights[2710];
				12'd2710	: data2 <= weights[2711];
				12'd2711	: data2 <= weights[2712];
				12'd2712	: data2 <= weights[2713];
				12'd2713	: data2 <= weights[2714];
				12'd2714	: data2 <= weights[2715];
				12'd2715	: data2 <= weights[2716];
				12'd2716	: data2 <= weights[2717];
				12'd2717	: data2 <= weights[2718];
				12'd2718	: data2 <= weights[2719];
				12'd2719	: data2 <= weights[2720];
				12'd2720	: data2 <= weights[2721];
				12'd2721	: data2 <= weights[2722];
				12'd2722	: data2 <= weights[2723];
				12'd2723	: data2 <= weights[2724];
				12'd2724	: data2 <= weights[2725];
				12'd2725	: data2 <= weights[2726];
				12'd2726	: data2 <= weights[2727];
				12'd2727	: data2 <= weights[2728];
				12'd2728	: data2 <= weights[2729];
				12'd2729	: data2 <= weights[2730];
				12'd2730	: data2 <= weights[2731];
				12'd2731	: data2 <= weights[2732];
				12'd2732	: data2 <= weights[2733];
				12'd2733	: data2 <= weights[2734];
				12'd2734	: data2 <= weights[2735];
				12'd2735	: data2 <= weights[2736];
				12'd2736	: data2 <= weights[2737];
				12'd2737	: data2 <= weights[2738];
				12'd2738	: data2 <= weights[2739];
				12'd2739	: data2 <= weights[2740];
				12'd2740	: data2 <= weights[2741];
				12'd2741	: data2 <= weights[2742];
				12'd2742	: data2 <= weights[2743];
				12'd2743	: data2 <= weights[2744];
				12'd2744	: data2 <= weights[2745];
				12'd2745	: data2 <= weights[2746];
				12'd2746	: data2 <= weights[2747];
				12'd2747	: data2 <= weights[2748];
				12'd2748	: data2 <= weights[2749];
				12'd2749	: data2 <= weights[2750];
				12'd2750	: data2 <= weights[2751];
				12'd2751	: data2 <= weights[2752];
				12'd2752	: data2 <= weights[2753];
				12'd2753	: data2 <= weights[2754];
				12'd2754	: data2 <= weights[2755];
				12'd2755	: data2 <= weights[2756];
				12'd2756	: data2 <= weights[2757];
				12'd2757	: data2 <= weights[2758];
				12'd2758	: data2 <= weights[2759];
				12'd2759	: data2 <= weights[2760];
				12'd2760	: data2 <= weights[2761];
				12'd2761	: data2 <= weights[2762];
				12'd2762	: data2 <= weights[2763];
				12'd2763	: data2 <= weights[2764];
				12'd2764	: data2 <= weights[2765];
				12'd2765	: data2 <= weights[2766];
				12'd2766	: data2 <= weights[2767];
				12'd2767	: data2 <= weights[2768];
				12'd2768	: data2 <= weights[2769];
				12'd2769	: data2 <= weights[2770];
				12'd2770	: data2 <= weights[2771];
				12'd2771	: data2 <= weights[2772];
				12'd2772	: data2 <= weights[2773];
				12'd2773	: data2 <= weights[2774];
				12'd2774	: data2 <= weights[2775];
				12'd2775	: data2 <= weights[2776];
				12'd2776	: data2 <= weights[2777];
				12'd2777	: data2 <= weights[2778];
				12'd2778	: data2 <= weights[2779];
				12'd2779	: data2 <= weights[2780];
				12'd2780	: data2 <= weights[2781];
				12'd2781	: data2 <= weights[2782];
				12'd2782	: data2 <= weights[2783];
				12'd2783	: data2 <= weights[2784];
				12'd2784	: data2 <= weights[2785];
				12'd2785	: data2 <= weights[2786];
				12'd2786	: data2 <= weights[2787];
				12'd2787	: data2 <= weights[2788];
				12'd2788	: data2 <= weights[2789];
				12'd2789	: data2 <= weights[2790];
				12'd2790	: data2 <= weights[2791];
				12'd2791	: data2 <= weights[2792];
				12'd2792	: data2 <= weights[2793];
				12'd2793	: data2 <= weights[2794];
				12'd2794	: data2 <= weights[2795];
				12'd2795	: data2 <= weights[2796];
				12'd2796	: data2 <= weights[2797];
				12'd2797	: data2 <= weights[2798];
				12'd2798	: data2 <= weights[2799];
				12'd2799	: data2 <= weights[2800];
				12'd2800	: data2 <= weights[2801];
				12'd2801	: data2 <= weights[2802];
				12'd2802	: data2 <= weights[2803];
				12'd2803	: data2 <= weights[2804];
				12'd2804	: data2 <= weights[2805];
				12'd2805	: data2 <= weights[2806];
				12'd2806	: data2 <= weights[2807];
				12'd2807	: data2 <= weights[2808];
				12'd2808	: data2 <= weights[2809];
				12'd2809	: data2 <= weights[2810];
				12'd2810	: data2 <= weights[2811];
				12'd2811	: data2 <= weights[2812];
				12'd2812	: data2 <= weights[2813];
				12'd2813	: data2 <= weights[2814];
				12'd2814	: data2 <= weights[2815];
				12'd2815	: data2 <= weights[2816];
				12'd2816	: data2 <= weights[2817];
				12'd2817	: data2 <= weights[2818];
				12'd2818	: data2 <= weights[2819];
				12'd2819	: data2 <= weights[2820];
				12'd2820	: data2 <= weights[2821];
				12'd2821	: data2 <= weights[2822];
				12'd2822	: data2 <= weights[2823];
				12'd2823	: data2 <= weights[2824];
				12'd2824	: data2 <= weights[2825];
				12'd2825	: data2 <= weights[2826];
				12'd2826	: data2 <= weights[2827];
				12'd2827	: data2 <= weights[2828];
				12'd2828	: data2 <= weights[2829];
				12'd2829	: data2 <= weights[2830];
				12'd2830	: data2 <= weights[2831];
				12'd2831	: data2 <= weights[2832];
				12'd2832	: data2 <= weights[2833];
				12'd2833	: data2 <= weights[2834];
				12'd2834	: data2 <= weights[2835];
				12'd2835	: data2 <= weights[2836];
				12'd2836	: data2 <= weights[2837];
				12'd2837	: data2 <= weights[2838];
				12'd2838	: data2 <= weights[2839];
				12'd2839	: data2 <= weights[2840];
				12'd2840	: data2 <= weights[2841];
				12'd2841	: data2 <= weights[2842];
				12'd2842	: data2 <= weights[2843];
				12'd2843	: data2 <= weights[2844];
				12'd2844	: data2 <= weights[2845];
				12'd2845	: data2 <= weights[2846];
				12'd2846	: data2 <= weights[2847];
				12'd2847	: data2 <= weights[2848];
				12'd2848	: data2 <= weights[2849];
				12'd2849	: data2 <= weights[2850];
				12'd2850	: data2 <= weights[2851];
				12'd2851	: data2 <= weights[2852];
				12'd2852	: data2 <= weights[2853];
				12'd2853	: data2 <= weights[2854];
				12'd2854	: data2 <= weights[2855];
				12'd2855	: data2 <= weights[2856];
				12'd2856	: data2 <= weights[2857];
				12'd2857	: data2 <= weights[2858];
				12'd2858	: data2 <= weights[2859];
				12'd2859	: data2 <= weights[2860];
				12'd2860	: data2 <= weights[2861];
				12'd2861	: data2 <= weights[2862];
				12'd2862	: data2 <= weights[2863];
				12'd2863	: data2 <= weights[2864];
				12'd2864	: data2 <= weights[2865];
				12'd2865	: data2 <= weights[2866];
				12'd2866	: data2 <= weights[2867];
				12'd2867	: data2 <= weights[2868];
				12'd2868	: data2 <= weights[2869];
				12'd2869	: data2 <= weights[2870];
				12'd2870	: data2 <= weights[2871];
				12'd2871	: data2 <= weights[2872];
				12'd2872	: data2 <= weights[2873];
				12'd2873	: data2 <= weights[2874];
				12'd2874	: data2 <= weights[2875];
				12'd2875	: data2 <= weights[2876];
				12'd2876	: data2 <= weights[2877];
				12'd2877	: data2 <= weights[2878];
				12'd2878	: data2 <= weights[2879];
				12'd2879	: data2 <= weights[2880];
				12'd2880	: data2 <= weights[2881];
				12'd2881	: data2 <= weights[2882];
				12'd2882	: data2 <= weights[2883];
				12'd2883	: data2 <= weights[2884];
				12'd2884	: data2 <= weights[2885];
				12'd2885	: data2 <= weights[2886];
				12'd2886	: data2 <= weights[2887];
				12'd2887	: data2 <= weights[2888];
				12'd2888	: data2 <= weights[2889];
				12'd2889	: data2 <= weights[2890];
				12'd2890	: data2 <= weights[2891];
				12'd2891	: data2 <= weights[2892];
				12'd2892	: data2 <= weights[2893];
				12'd2893	: data2 <= weights[2894];
				12'd2894	: data2 <= weights[2895];
				12'd2895	: data2 <= weights[2896];
				12'd2896	: data2 <= weights[2897];
				12'd2897	: data2 <= weights[2898];
				12'd2898	: data2 <= weights[2899];
				12'd2899	: data2 <= weights[2900];
				12'd2900	: data2 <= weights[2901];
				12'd2901	: data2 <= weights[2902];
				12'd2902	: data2 <= weights[2903];
				12'd2903	: data2 <= weights[2904];
				12'd2904	: data2 <= weights[2905];
				12'd2905	: data2 <= weights[2906];
				12'd2906	: data2 <= weights[2907];
				12'd2907	: data2 <= weights[2908];
				12'd2908	: data2 <= weights[2909];
				12'd2909	: data2 <= weights[2910];
				12'd2910	: data2 <= weights[2911];
				12'd2911	: data2 <= weights[2912];
				12'd2912	: data2 <= weights[2913];
				12'd2913	: data2 <= weights[2914];
				12'd2914	: data2 <= weights[2915];
				12'd2915	: data2 <= weights[2916];
				12'd2916	: data2 <= weights[2917];
				12'd2917	: data2 <= weights[2918];
				12'd2918	: data2 <= weights[2919];
				12'd2919	: data2 <= weights[2920];
				12'd2920	: data2 <= weights[2921];
				12'd2921	: data2 <= weights[2922];
				12'd2922	: data2 <= weights[2923];
				12'd2923	: data2 <= weights[2924];
				12'd2924	: data2 <= weights[2925];
				12'd2925	: data2 <= weights[2926];
				12'd2926	: data2 <= weights[2927];
				12'd2927	: data2 <= weights[2928];
				12'd2928	: data2 <= weights[2929];
				12'd2929	: data2 <= weights[2930];
				12'd2930	: data2 <= weights[2931];
				12'd2931	: data2 <= weights[2932];
				12'd2932	: data2 <= weights[2933];
				12'd2933	: data2 <= weights[2934];
				12'd2934	: data2 <= weights[2935];
				12'd2935	: data2 <= weights[2936];
				12'd2936	: data2 <= weights[2937];
				12'd2937	: data2 <= weights[2938];
				12'd2938	: data2 <= weights[2939];
				12'd2939	: data2 <= weights[2940];
				12'd2940	: data2 <= weights[2941];
				12'd2941	: data2 <= weights[2942];
				12'd2942	: data2 <= weights[2943];
				12'd2943	: data2 <= weights[2944];
				12'd2944	: data2 <= weights[2945];
				12'd2945	: data2 <= weights[2946];
				12'd2946	: data2 <= weights[2947];
				12'd2947	: data2 <= weights[2948];
				12'd2948	: data2 <= weights[2949];
				12'd2949	: data2 <= weights[2950];
				12'd2950	: data2 <= weights[2951];
				12'd2951	: data2 <= weights[2952];
				12'd2952	: data2 <= weights[2953];
				12'd2953	: data2 <= weights[2954];
				12'd2954	: data2 <= weights[2955];
				12'd2955	: data2 <= weights[2956];
				12'd2956	: data2 <= weights[2957];
				12'd2957	: data2 <= weights[2958];
				12'd2958	: data2 <= weights[2959];
				12'd2959	: data2 <= weights[2960];
				12'd2960	: data2 <= weights[2961];
				12'd2961	: data2 <= weights[2962];
				12'd2962	: data2 <= weights[2963];
				12'd2963	: data2 <= weights[2964];
				12'd2964	: data2 <= weights[2965];
				12'd2965	: data2 <= weights[2966];
				12'd2966	: data2 <= weights[2967];
				12'd2967	: data2 <= weights[2968];
				12'd2968	: data2 <= weights[2969];
				12'd2969	: data2 <= weights[2970];
				12'd2970	: data2 <= weights[2971];
				12'd2971	: data2 <= weights[2972];
				12'd2972	: data2 <= weights[2973];
				12'd2973	: data2 <= weights[2974];
				12'd2974	: data2 <= weights[2975];
				12'd2975	: data2 <= weights[2976];
				12'd2976	: data2 <= weights[2977];
				12'd2977	: data2 <= weights[2978];
				12'd2978	: data2 <= weights[2979];
				12'd2979	: data2 <= weights[2980];
				12'd2980	: data2 <= weights[2981];
				12'd2981	: data2 <= weights[2982];
				12'd2982	: data2 <= weights[2983];
				12'd2983	: data2 <= weights[2984];
				12'd2984	: data2 <= weights[2985];
				12'd2985	: data2 <= weights[2986];
				12'd2986	: data2 <= weights[2987];
				12'd2987	: data2 <= weights[2988];
				12'd2988	: data2 <= weights[2989];
				12'd2989	: data2 <= weights[2990];
				12'd2990	: data2 <= weights[2991];
				12'd2991	: data2 <= weights[2992];
				12'd2992	: data2 <= weights[2993];
				12'd2993	: data2 <= weights[2994];
				12'd2994	: data2 <= weights[2995];
				12'd2995	: data2 <= weights[2996];
				12'd2996	: data2 <= weights[2997];
				12'd2997	: data2 <= weights[2998];
				12'd2998	: data2 <= weights[2999];
				12'd2999	: data2 <= weights[3000];
				12'd3000	: data2 <= weights[3001];
				12'd3001	: data2 <= weights[3002];
				12'd3002	: data2 <= weights[3003];
				12'd3003	: data2 <= weights[3004];
				12'd3004	: data2 <= weights[3005];
				12'd3005	: data2 <= weights[3006];
				12'd3006	: data2 <= weights[3007];
				12'd3007	: data2 <= weights[3008];
				12'd3008	: data2 <= weights[3009];
				12'd3009	: data2 <= weights[3010];
				12'd3010	: data2 <= weights[3011];
				12'd3011	: data2 <= weights[3012];
				12'd3012	: data2 <= weights[3013];
				12'd3013	: data2 <= weights[3014];
				12'd3014	: data2 <= weights[3015];
				12'd3015	: data2 <= weights[3016];
				12'd3016	: data2 <= weights[3017];
				12'd3017	: data2 <= weights[3018];
				12'd3018	: data2 <= weights[3019];
				12'd3019	: data2 <= weights[3020];
				12'd3020	: data2 <= weights[3021];
				12'd3021	: data2 <= weights[3022];
				12'd3022	: data2 <= weights[3023];
				12'd3023	: data2 <= weights[3024];
				12'd3024	: data2 <= weights[3025];
				12'd3025	: data2 <= weights[3026];
				12'd3026	: data2 <= weights[3027];
				12'd3027	: data2 <= weights[3028];
				12'd3028	: data2 <= weights[3029];
				12'd3029	: data2 <= weights[3030];
				12'd3030	: data2 <= weights[3031];
				12'd3031	: data2 <= weights[3032];
				12'd3032	: data2 <= weights[3033];
				12'd3033	: data2 <= weights[3034];
				12'd3034	: data2 <= weights[3035];
				12'd3035	: data2 <= weights[3036];
				12'd3036	: data2 <= weights[3037];
				12'd3037	: data2 <= weights[3038];
				12'd3038	: data2 <= weights[3039];
				12'd3039	: data2 <= weights[3040];
				12'd3040	: data2 <= weights[3041];
				12'd3041	: data2 <= weights[3042];
				12'd3042	: data2 <= weights[3043];
				12'd3043	: data2 <= weights[3044];
				12'd3044	: data2 <= weights[3045];
				12'd3045	: data2 <= weights[3046];
				12'd3046	: data2 <= weights[3047];
				12'd3047	: data2 <= weights[3048];
				12'd3048	: data2 <= weights[3049];
				12'd3049	: data2 <= weights[3050];
				12'd3050	: data2 <= weights[3051];
				12'd3051	: data2 <= weights[3052];
				12'd3052	: data2 <= weights[3053];
				12'd3053	: data2 <= weights[3054];
				12'd3054	: data2 <= weights[3055];
				12'd3055	: data2 <= weights[3056];
				12'd3056	: data2 <= weights[3057];
				12'd3057	: data2 <= weights[3058];
				12'd3058	: data2 <= weights[3059];
				12'd3059	: data2 <= weights[3060];
				12'd3060	: data2 <= weights[3061];
				12'd3061	: data2 <= weights[3062];
				12'd3062	: data2 <= weights[3063];
				12'd3063	: data2 <= weights[3064];
				12'd3064	: data2 <= weights[3065];
				12'd3065	: data2 <= weights[3066];
				12'd3066	: data2 <= weights[3067];
				12'd3067	: data2 <= weights[3068];
				12'd3068	: data2 <= weights[3069];
				12'd3069	: data2 <= weights[3070];
				12'd3070	: data2 <= weights[3071];
				12'd3071	: data2 <= weights[3072];
				12'd3072	: data2 <= weights[3073];
				12'd3073	: data2 <= weights[3074];
				12'd3074	: data2 <= weights[3075];
				12'd3075	: data2 <= weights[3076];
				12'd3076	: data2 <= weights[3077];
				12'd3077	: data2 <= weights[3078];
				12'd3078	: data2 <= weights[3079];
				12'd3079	: data2 <= weights[3080];
				12'd3080	: data2 <= weights[3081];
				12'd3081	: data2 <= weights[3082];
				12'd3082	: data2 <= weights[3083];
				12'd3083	: data2 <= weights[3084];
				12'd3084	: data2 <= weights[3085];
				12'd3085	: data2 <= weights[3086];
				12'd3086	: data2 <= weights[3087];
				12'd3087	: data2 <= weights[3088];
				12'd3088	: data2 <= weights[3089];
				12'd3089	: data2 <= weights[3090];
				12'd3090	: data2 <= weights[3091];
				12'd3091	: data2 <= weights[3092];
				12'd3092	: data2 <= weights[3093];
				12'd3093	: data2 <= weights[3094];
				12'd3094	: data2 <= weights[3095];
				12'd3095	: data2 <= weights[3096];
				12'd3096	: data2 <= weights[3097];
				12'd3097	: data2 <= weights[3098];
				12'd3098	: data2 <= weights[3099];
				12'd3099	: data2 <= weights[3100];
				12'd3100	: data2 <= weights[3101];
				12'd3101	: data2 <= weights[3102];
				12'd3102	: data2 <= weights[3103];
				12'd3103	: data2 <= weights[3104];
				12'd3104	: data2 <= weights[3105];
				12'd3105	: data2 <= weights[3106];
				12'd3106	: data2 <= weights[3107];
				12'd3107	: data2 <= weights[3108];
				12'd3108	: data2 <= weights[3109];
				12'd3109	: data2 <= weights[3110];
				12'd3110	: data2 <= weights[3111];
				12'd3111	: data2 <= weights[3112];
				12'd3112	: data2 <= weights[3113];
				12'd3113	: data2 <= weights[3114];
				12'd3114	: data2 <= weights[3115];
				12'd3115	: data2 <= weights[3116];
				12'd3116	: data2 <= weights[3117];
				12'd3117	: data2 <= weights[3118];
				12'd3118	: data2 <= weights[3119];
				12'd3119	: data2 <= weights[3120];
				12'd3120	: data2 <= weights[3121];
				12'd3121	: data2 <= weights[3122];
				12'd3122	: data2 <= weights[3123];
				12'd3123	: data2 <= weights[3124];
				12'd3124	: data2 <= weights[3125];
				12'd3125	: data2 <= weights[3126];
				12'd3126	: data2 <= weights[3127];
				12'd3127	: data2 <= weights[3128];
				12'd3128	: data2 <= weights[3129];
				12'd3129	: data2 <= weights[3130];
				12'd3130	: data2 <= weights[3131];
				12'd3131	: data2 <= weights[3132];
				12'd3132	: data2 <= weights[3133];
				12'd3133	: data2 <= weights[3134];
				12'd3134	: data2 <= weights[3135];
				12'd3135	: data2 <= weights[3136];
				12'd3136	: data2 <= weights[3137];
				12'd3137	: data2 <= weights[3138];
				12'd3138	: data2 <= weights[3139];
				12'd3139	: data2 <= weights[3140];
				12'd3140	: data2 <= weights[3141];
				12'd3141	: data2 <= weights[3142];
				12'd3142	: data2 <= weights[3143];
				12'd3143	: data2 <= weights[3144];
				12'd3144	: data2 <= weights[3145];
				12'd3145	: data2 <= weights[3146];
				12'd3146	: data2 <= weights[3147];
				12'd3147	: data2 <= weights[3148];
				12'd3148	: data2 <= weights[3149];
				12'd3149	: data2 <= weights[3150];
				12'd3150	: data2 <= weights[3151];
				12'd3151	: data2 <= weights[3152];
				12'd3152	: data2 <= weights[3153];
				12'd3153	: data2 <= weights[3154];
				12'd3154	: data2 <= weights[3155];
				12'd3155	: data2 <= weights[3156];
				12'd3156	: data2 <= weights[3157];
				12'd3157	: data2 <= weights[3158];
				12'd3158	: data2 <= weights[3159];
				12'd3159	: data2 <= weights[3160];
				12'd3160	: data2 <= weights[3161];
				12'd3161	: data2 <= weights[3162];
				12'd3162	: data2 <= weights[3163];
				12'd3163	: data2 <= weights[3164];
				12'd3164	: data2 <= weights[3165];
				12'd3165	: data2 <= weights[3166];
				12'd3166	: data2 <= weights[3167];
				12'd3167	: data2 <= weights[3168];
				12'd3168	: data2 <= weights[3169];
				12'd3169	: data2 <= weights[3170];
				12'd3170	: data2 <= weights[3171];
				12'd3171	: data2 <= weights[3172];
				12'd3172	: data2 <= weights[3173];
				12'd3173	: data2 <= weights[3174];
				12'd3174	: data2 <= weights[3175];
				12'd3175	: data2 <= weights[3176];
				12'd3176	: data2 <= weights[3177];
				12'd3177	: data2 <= weights[3178];
				12'd3178	: data2 <= weights[3179];
				12'd3179	: data2 <= weights[3180];
				12'd3180	: data2 <= weights[3181];
				12'd3181	: data2 <= weights[3182];
				12'd3182	: data2 <= weights[3183];
				12'd3183	: data2 <= weights[3184];
				12'd3184	: data2 <= weights[3185];
				12'd3185	: data2 <= weights[3186];
				12'd3186	: data2 <= weights[3187];
				12'd3187	: data2 <= weights[3188];
				12'd3188	: data2 <= weights[3189];
				12'd3189	: data2 <= weights[3190];
				12'd3190	: data2 <= weights[3191];
				12'd3191	: data2 <= weights[3192];
				12'd3192	: data2 <= weights[3193];
				12'd3193	: data2 <= weights[3194];
				12'd3194	: data2 <= weights[3195];
				12'd3195	: data2 <= weights[3196];
				12'd3196	: data2 <= weights[3197];
				12'd3197	: data2 <= weights[3198];
				12'd3198	: data2 <= weights[3199];
				12'd3199	: data2 <= weights[3200];
				12'd3200	: data2 <= weights[3201];
				12'd3201	: data2 <= weights[3202];
				12'd3202	: data2 <= weights[3203];
				12'd3203	: data2 <= weights[3204];
				12'd3204	: data2 <= weights[3205];
				12'd3205	: data2 <= weights[3206];
				12'd3206	: data2 <= weights[3207];
				12'd3207	: data2 <= weights[3208];
				12'd3208	: data2 <= weights[3209];
				12'd3209	: data2 <= weights[3210];
				12'd3210	: data2 <= weights[3211];
				12'd3211	: data2 <= weights[3212];
				12'd3212	: data2 <= weights[3213];
				12'd3213	: data2 <= weights[3214];
				12'd3214	: data2 <= weights[3215];
				12'd3215	: data2 <= weights[3216];
				12'd3216	: data2 <= weights[3217];
				12'd3217	: data2 <= weights[3218];
				12'd3218	: data2 <= weights[3219];
				12'd3219	: data2 <= weights[3220];
				12'd3220	: data2 <= weights[3221];
				12'd3221	: data2 <= weights[3222];
				12'd3222	: data2 <= weights[3223];
				12'd3223	: data2 <= weights[3224];
				12'd3224	: data2 <= weights[3225];
				12'd3225	: data2 <= weights[3226];
				12'd3226	: data2 <= weights[3227];
				12'd3227	: data2 <= weights[3228];
				12'd3228	: data2 <= weights[3229];
				12'd3229	: data2 <= weights[3230];
				12'd3230	: data2 <= weights[3231];
				12'd3231	: data2 <= weights[3232];
				12'd3232	: data2 <= weights[3233];
				12'd3233	: data2 <= weights[3234];
				12'd3234	: data2 <= weights[3235];
				12'd3235	: data2 <= weights[3236];
				12'd3236	: data2 <= weights[3237];
				12'd3237	: data2 <= weights[3238];
				12'd3238	: data2 <= weights[3239];
				12'd3239	: data2 <= weights[3240];
				12'd3240	: data2 <= weights[3241];
				12'd3241	: data2 <= weights[3242];
				12'd3242	: data2 <= weights[3243];
				12'd3243	: data2 <= weights[3244];
				12'd3244	: data2 <= weights[3245];
				12'd3245	: data2 <= weights[3246];
				12'd3246	: data2 <= weights[3247];
				12'd3247	: data2 <= weights[3248];
				12'd3248	: data2 <= weights[3249];
				12'd3249	: data2 <= weights[3250];
				12'd3250	: data2 <= weights[3251];
				12'd3251	: data2 <= weights[3252];
				12'd3252	: data2 <= weights[3253];
				12'd3253	: data2 <= weights[3254];
				12'd3254	: data2 <= weights[3255];
				12'd3255	: data2 <= weights[3256];
				12'd3256	: data2 <= weights[3257];
				12'd3257	: data2 <= weights[3258];
				12'd3258	: data2 <= weights[3259];
				12'd3259	: data2 <= weights[3260];
				12'd3260	: data2 <= weights[3261];
				12'd3261	: data2 <= weights[3262];
				12'd3262	: data2 <= weights[3263];
				12'd3263	: data2 <= weights[3264];
				12'd3264	: data2 <= weights[3265];
				12'd3265	: data2 <= weights[3266];
				12'd3266	: data2 <= weights[3267];
				12'd3267	: data2 <= weights[3268];
				12'd3268	: data2 <= weights[3269];
				12'd3269	: data2 <= weights[3270];
				12'd3270	: data2 <= weights[3271];
				12'd3271	: data2 <= weights[3272];
				12'd3272	: data2 <= weights[3273];
				12'd3273	: data2 <= weights[3274];
				12'd3274	: data2 <= weights[3275];
				12'd3275	: data2 <= weights[3276];
				12'd3276	: data2 <= weights[3277];
				12'd3277	: data2 <= weights[3278];
				12'd3278	: data2 <= weights[3279];
				12'd3279	: data2 <= weights[3280];
				12'd3280	: data2 <= weights[3281];
				12'd3281	: data2 <= weights[3282];
				12'd3282	: data2 <= weights[3283];
				12'd3283	: data2 <= weights[3284];
				12'd3284	: data2 <= weights[3285];
				12'd3285	: data2 <= weights[3286];
				12'd3286	: data2 <= weights[3287];
				12'd3287	: data2 <= weights[3288];
				12'd3288	: data2 <= weights[3289];
				12'd3289	: data2 <= weights[3290];
				12'd3290	: data2 <= weights[3291];
				12'd3291	: data2 <= weights[3292];
				12'd3292	: data2 <= weights[3293];
				12'd3293	: data2 <= weights[3294];
				12'd3294	: data2 <= weights[3295];
				12'd3295	: data2 <= weights[3296];
				12'd3296	: data2 <= weights[3297];
				12'd3297	: data2 <= weights[3298];
				12'd3298	: data2 <= weights[3299];
				12'd3299	: data2 <= weights[3300];
				12'd3300	: data2 <= weights[3301];
				12'd3301	: data2 <= weights[3302];
				12'd3302	: data2 <= weights[3303];
				12'd3303	: data2 <= weights[3304];
				12'd3304	: data2 <= weights[3305];
				12'd3305	: data2 <= weights[3306];
				12'd3306	: data2 <= weights[3307];
				12'd3307	: data2 <= weights[3308];
				12'd3308	: data2 <= weights[3309];
				12'd3309	: data2 <= weights[3310];
				12'd3310	: data2 <= weights[3311];
				12'd3311	: data2 <= weights[3312];
				12'd3312	: data2 <= weights[3313];
				12'd3313	: data2 <= weights[3314];
				12'd3314	: data2 <= weights[3315];
				12'd3315	: data2 <= weights[3316];
				12'd3316	: data2 <= weights[3317];
				12'd3317	: data2 <= weights[3318];
				12'd3318	: data2 <= weights[3319];
				12'd3319	: data2 <= weights[3320];
				12'd3320	: data2 <= weights[3321];
				12'd3321	: data2 <= weights[3322];
				12'd3322	: data2 <= weights[3323];
				12'd3323	: data2 <= weights[3324];
				12'd3324	: data2 <= weights[3325];
				12'd3325	: data2 <= weights[3326];
				12'd3326	: data2 <= weights[3327];
				12'd3327	: data2 <= weights[3328];
				12'd3328	: data2 <= weights[3329];
				12'd3329	: data2 <= weights[3330];
				12'd3330	: data2 <= weights[3331];
				12'd3331	: data2 <= weights[3332];
				12'd3332	: data2 <= weights[3333];
				12'd3333	: data2 <= weights[3334];
				12'd3334	: data2 <= weights[3335];
				12'd3335	: data2 <= weights[3336];
				12'd3336	: data2 <= weights[3337];
				12'd3337	: data2 <= weights[3338];
				12'd3338	: data2 <= weights[3339];
				12'd3339	: data2 <= weights[3340];
				12'd3340	: data2 <= weights[3341];
				12'd3341	: data2 <= weights[3342];
				12'd3342	: data2 <= weights[3343];
				12'd3343	: data2 <= weights[3344];
				12'd3344	: data2 <= weights[3345];
				12'd3345	: data2 <= weights[3346];
				12'd3346	: data2 <= weights[3347];
				12'd3347	: data2 <= weights[3348];
				12'd3348	: data2 <= weights[3349];
				12'd3349	: data2 <= weights[3350];
				12'd3350	: data2 <= weights[3351];
				12'd3351	: data2 <= weights[3352];
				12'd3352	: data2 <= weights[3353];
				12'd3353	: data2 <= weights[3354];
				12'd3354	: data2 <= weights[3355];
				12'd3355	: data2 <= weights[3356];
				12'd3356	: data2 <= weights[3357];
				12'd3357	: data2 <= weights[3358];
				12'd3358	: data2 <= weights[3359];
				12'd3359	: data2 <= weights[3360];
				12'd3360	: data2 <= weights[3361];
				12'd3361	: data2 <= weights[3362];
				12'd3362	: data2 <= weights[3363];
				12'd3363	: data2 <= weights[3364];
				12'd3364	: data2 <= weights[3365];
				12'd3365	: data2 <= weights[3366];
				12'd3366	: data2 <= weights[3367];
				12'd3367	: data2 <= weights[3368];
				12'd3368	: data2 <= weights[3369];
				12'd3369	: data2 <= weights[3370];
				12'd3370	: data2 <= weights[3371];
				12'd3371	: data2 <= weights[3372];
				12'd3372	: data2 <= weights[3373];
				12'd3373	: data2 <= weights[3374];
				12'd3374	: data2 <= weights[3375];
				12'd3375	: data2 <= weights[3376];
				12'd3376	: data2 <= weights[3377];
				12'd3377	: data2 <= weights[3378];
				12'd3378	: data2 <= weights[3379];
				12'd3379	: data2 <= weights[3380];
				12'd3380	: data2 <= weights[3381];
				12'd3381	: data2 <= weights[3382];
				12'd3382	: data2 <= weights[3383];
				12'd3383	: data2 <= weights[3384];
				12'd3384	: data2 <= weights[3385];
				12'd3385	: data2 <= weights[3386];
				12'd3386	: data2 <= weights[3387];
				12'd3387	: data2 <= weights[3388];
				12'd3388	: data2 <= weights[3389];
				12'd3389	: data2 <= weights[3390];
				12'd3390	: data2 <= weights[3391];
				12'd3391	: data2 <= weights[3392];
				12'd3392	: data2 <= weights[3393];
				12'd3393	: data2 <= weights[3394];
				12'd3394	: data2 <= weights[3395];
				12'd3395	: data2 <= weights[3396];
				12'd3396	: data2 <= weights[3397];
				12'd3397	: data2 <= weights[3398];
				12'd3398	: data2 <= weights[3399];
				12'd3399	: data2 <= weights[3400];
				12'd3400	: data2 <= weights[3401];
				12'd3401	: data2 <= weights[3402];
				12'd3402	: data2 <= weights[3403];
				12'd3403	: data2 <= weights[3404];
				12'd3404	: data2 <= weights[3405];
				12'd3405	: data2 <= weights[3406];
				12'd3406	: data2 <= weights[3407];
				12'd3407	: data2 <= weights[3408];
				12'd3408	: data2 <= weights[3409];
				12'd3409	: data2 <= weights[3410];
				12'd3410	: data2 <= weights[3411];
				12'd3411	: data2 <= weights[3412];
				12'd3412	: data2 <= weights[3413];
				12'd3413	: data2 <= weights[3414];
				12'd3414	: data2 <= weights[3415];
				12'd3415	: data2 <= weights[3416];
				12'd3416	: data2 <= weights[3417];
				12'd3417	: data2 <= weights[3418];
				12'd3418	: data2 <= weights[3419];
				12'd3419	: data2 <= weights[3420];
				12'd3420	: data2 <= weights[3421];
				12'd3421	: data2 <= weights[3422];
				12'd3422	: data2 <= weights[3423];
				12'd3423	: data2 <= weights[3424];
				12'd3424	: data2 <= weights[3425];
				12'd3425	: data2 <= weights[3426];
				12'd3426	: data2 <= weights[3427];
				12'd3427	: data2 <= weights[3428];
				12'd3428	: data2 <= weights[3429];
				12'd3429	: data2 <= weights[3430];
				12'd3430	: data2 <= weights[3431];
				12'd3431	: data2 <= weights[3432];
				12'd3432	: data2 <= weights[3433];
				12'd3433	: data2 <= weights[3434];
				12'd3434	: data2 <= weights[3435];
				12'd3435	: data2 <= weights[3436];
				12'd3436	: data2 <= weights[3437];
				12'd3437	: data2 <= weights[3438];
				12'd3438	: data2 <= weights[3439];
				12'd3439	: data2 <= weights[3440];
				12'd3440	: data2 <= weights[3441];
				12'd3441	: data2 <= weights[3442];
				12'd3442	: data2 <= weights[3443];
				12'd3443	: data2 <= weights[3444];
				12'd3444	: data2 <= weights[3445];
				12'd3445	: data2 <= weights[3446];
				12'd3446	: data2 <= weights[3447];
				12'd3447	: data2 <= weights[3448];
				12'd3448	: data2 <= weights[3449];
				12'd3449	: data2 <= weights[3450];
				12'd3450	: data2 <= weights[3451];
				12'd3451	: data2 <= weights[3452];
				12'd3452	: data2 <= weights[3453];
				12'd3453	: data2 <= weights[3454];
				12'd3454	: data2 <= weights[3455];
				12'd3455	: data2 <= weights[3456];
				12'd3456	: data2 <= weights[3457];
				12'd3457	: data2 <= weights[3458];
				12'd3458	: data2 <= weights[3459];
				12'd3459	: data2 <= weights[3460];
				12'd3460	: data2 <= weights[3461];
				12'd3461	: data2 <= weights[3462];
				12'd3462	: data2 <= weights[3463];
				12'd3463	: data2 <= weights[3464];
				12'd3464	: data2 <= weights[3465];
				12'd3465	: data2 <= weights[3466];
				12'd3466	: data2 <= weights[3467];
				12'd3467	: data2 <= weights[3468];
				12'd3468	: data2 <= weights[3469];
				12'd3469	: data2 <= weights[3470];
				12'd3470	: data2 <= weights[3471];
				12'd3471	: data2 <= weights[3472];
				12'd3472	: data2 <= weights[3473];
				12'd3473	: data2 <= weights[3474];
				12'd3474	: data2 <= weights[3475];
				12'd3475	: data2 <= weights[3476];
				12'd3476	: data2 <= weights[3477];
				12'd3477	: data2 <= weights[3478];
				12'd3478	: data2 <= weights[3479];
				12'd3479	: data2 <= weights[3480];
				12'd3480	: data2 <= weights[3481];
				12'd3481	: data2 <= weights[3482];
				12'd3482	: data2 <= weights[3483];
				12'd3483	: data2 <= weights[3484];
				12'd3484	: data2 <= weights[3485];
				12'd3485	: data2 <= weights[3486];
				12'd3486	: data2 <= weights[3487];
				12'd3487	: data2 <= weights[3488];
				12'd3488	: data2 <= weights[3489];
				12'd3489	: data2 <= weights[3490];
				12'd3490	: data2 <= weights[3491];
				12'd3491	: data2 <= weights[3492];
				12'd3492	: data2 <= weights[3493];
				12'd3493	: data2 <= weights[3494];
				12'd3494	: data2 <= weights[3495];
				12'd3495	: data2 <= weights[3496];
				12'd3496	: data2 <= weights[3497];
				12'd3497	: data2 <= weights[3498];
				12'd3498	: data2 <= weights[3499];
				12'd3499	: data2 <= weights[3500];
				12'd3500	: data2 <= weights[3501];
				12'd3501	: data2 <= weights[3502];
				12'd3502	: data2 <= weights[3503];
				12'd3503	: data2 <= weights[3504];
				12'd3504	: data2 <= weights[3505];
				12'd3505	: data2 <= weights[3506];
				12'd3506	: data2 <= weights[3507];
				12'd3507	: data2 <= weights[3508];
				12'd3508	: data2 <= weights[3509];
				12'd3509	: data2 <= weights[3510];
				12'd3510	: data2 <= weights[3511];
				12'd3511	: data2 <= weights[3512];
				12'd3512	: data2 <= weights[3513];
				12'd3513	: data2 <= weights[3514];
				12'd3514	: data2 <= weights[3515];
				12'd3515	: data2 <= weights[3516];
				12'd3516	: data2 <= weights[3517];
				12'd3517	: data2 <= weights[3518];
				12'd3518	: data2 <= weights[3519];
				12'd3519	: data2 <= weights[3520];
				12'd3520	: data2 <= weights[3521];
				12'd3521	: data2 <= weights[3522];
				12'd3522	: data2 <= weights[3523];
				12'd3523	: data2 <= weights[3524];
				12'd3524	: data2 <= weights[3525];
				12'd3525	: data2 <= weights[3526];
				12'd3526	: data2 <= weights[3527];
				12'd3527	: data2 <= weights[3528];
				12'd3528	: data2 <= weights[3529];
				12'd3529	: data2 <= weights[3530];
				12'd3530	: data2 <= weights[3531];
				12'd3531	: data2 <= weights[3532];
				12'd3532	: data2 <= weights[3533];
				12'd3533	: data2 <= weights[3534];
				12'd3534	: data2 <= weights[3535];
				12'd3535	: data2 <= weights[3536];
				12'd3536	: data2 <= weights[3537];
				12'd3537	: data2 <= weights[3538];
				12'd3538	: data2 <= weights[3539];
				12'd3539	: data2 <= weights[3540];
				12'd3540	: data2 <= weights[3541];
				12'd3541	: data2 <= weights[3542];
				12'd3542	: data2 <= weights[3543];
				12'd3543	: data2 <= weights[3544];
				12'd3544	: data2 <= weights[3545];
				12'd3545	: data2 <= weights[3546];
				12'd3546	: data2 <= weights[3547];
				12'd3547	: data2 <= weights[3548];
				12'd3548	: data2 <= weights[3549];
				12'd3549	: data2 <= weights[3550];
				12'd3550	: data2 <= weights[3551];
				12'd3551	: data2 <= weights[3552];
				12'd3552	: data2 <= weights[3553];
				12'd3553	: data2 <= weights[3554];
				12'd3554	: data2 <= weights[3555];
				12'd3555	: data2 <= weights[3556];
				12'd3556	: data2 <= weights[3557];
				12'd3557	: data2 <= weights[3558];
				12'd3558	: data2 <= weights[3559];
				12'd3559	: data2 <= weights[3560];
				12'd3560	: data2 <= weights[3561];
				12'd3561	: data2 <= weights[3562];
				12'd3562	: data2 <= weights[3563];
				12'd3563	: data2 <= weights[3564];
				12'd3564	: data2 <= weights[3565];
				12'd3565	: data2 <= weights[3566];
				12'd3566	: data2 <= weights[3567];
				12'd3567	: data2 <= weights[3568];
				12'd3568	: data2 <= weights[3569];
				12'd3569	: data2 <= weights[3570];
				12'd3570	: data2 <= weights[3571];
				12'd3571	: data2 <= weights[3572];
				12'd3572	: data2 <= weights[3573];
				12'd3573	: data2 <= weights[3574];
				12'd3574	: data2 <= weights[3575];
				12'd3575	: data2 <= weights[3576];
				12'd3576	: data2 <= weights[3577];
				12'd3577	: data2 <= weights[3578];
				12'd3578	: data2 <= weights[3579];
				12'd3579	: data2 <= weights[3580];
				12'd3580	: data2 <= weights[3581];
				12'd3581	: data2 <= weights[3582];
				12'd3582	: data2 <= weights[3583];
				12'd3583	: data2 <= weights[3584];
				12'd3584	: data2 <= weights[3585];
				12'd3585	: data2 <= weights[3586];
				12'd3586	: data2 <= weights[3587];
				12'd3587	: data2 <= weights[3588];
				12'd3588	: data2 <= weights[3589];
				12'd3589	: data2 <= weights[3590];
				12'd3590	: data2 <= weights[3591];
				12'd3591	: data2 <= weights[3592];
				12'd3592	: data2 <= weights[3593];
				12'd3593	: data2 <= weights[3594];
				12'd3594	: data2 <= weights[3595];
				12'd3595	: data2 <= weights[3596];
				12'd3596	: data2 <= weights[3597];
				12'd3597	: data2 <= weights[3598];
				12'd3598	: data2 <= weights[3599];
				12'd3599	: data2 <= weights[3600];
				12'd3600	: data2 <= weights[3601];
				12'd3601	: data2 <= weights[3602];
				12'd3602	: data2 <= weights[3603];
				12'd3603	: data2 <= weights[3604];
				12'd3604	: data2 <= weights[3605];
				12'd3605	: data2 <= weights[3606];
				12'd3606	: data2 <= weights[3607];
				12'd3607	: data2 <= weights[3608];
				12'd3608	: data2 <= weights[3609];
				12'd3609	: data2 <= weights[3610];
				12'd3610	: data2 <= weights[3611];
				12'd3611	: data2 <= weights[3612];
				12'd3612	: data2 <= weights[3613];
				12'd3613	: data2 <= weights[3614];
				12'd3614	: data2 <= weights[3615];
				12'd3615	: data2 <= weights[3616];
				12'd3616	: data2 <= weights[3617];
				12'd3617	: data2 <= weights[3618];
				12'd3618	: data2 <= weights[3619];
				12'd3619	: data2 <= weights[3620];
				12'd3620	: data2 <= weights[3621];
				12'd3621	: data2 <= weights[3622];
				12'd3622	: data2 <= weights[3623];
				12'd3623	: data2 <= weights[3624];
				12'd3624	: data2 <= weights[3625];
				12'd3625	: data2 <= weights[3626];
				12'd3626	: data2 <= weights[3627];
				12'd3627	: data2 <= weights[3628];
				12'd3628	: data2 <= weights[3629];
				12'd3629	: data2 <= weights[3630];
				12'd3630	: data2 <= weights[3631];
				12'd3631	: data2 <= weights[3632];
				12'd3632	: data2 <= weights[3633];
				12'd3633	: data2 <= weights[3634];
				12'd3634	: data2 <= weights[3635];
				12'd3635	: data2 <= weights[3636];
				12'd3636	: data2 <= weights[3637];
				12'd3637	: data2 <= weights[3638];
				12'd3638	: data2 <= weights[3639];
				12'd3639	: data2 <= weights[3640];
				12'd3640	: data2 <= weights[3641];
				12'd3641	: data2 <= weights[3642];
				12'd3642	: data2 <= weights[3643];
				12'd3643	: data2 <= weights[3644];
				12'd3644	: data2 <= weights[3645];
				12'd3645	: data2 <= weights[3646];
				12'd3646	: data2 <= weights[3647];
				12'd3647	: data2 <= weights[3648];
				12'd3648	: data2 <= weights[3649];
				12'd3649	: data2 <= weights[3650];
				12'd3650	: data2 <= weights[3651];
				12'd3651	: data2 <= weights[3652];
				12'd3652	: data2 <= weights[3653];
				12'd3653	: data2 <= weights[3654];
				12'd3654	: data2 <= weights[3655];
				12'd3655	: data2 <= weights[3656];
				12'd3656	: data2 <= weights[3657];
				12'd3657	: data2 <= weights[3658];
				12'd3658	: data2 <= weights[3659];
				12'd3659	: data2 <= weights[3660];
				12'd3660	: data2 <= weights[3661];
				12'd3661	: data2 <= weights[3662];
				12'd3662	: data2 <= weights[3663];
				12'd3663	: data2 <= weights[3664];
				12'd3664	: data2 <= weights[3665];
				12'd3665	: data2 <= weights[3666];
				12'd3666	: data2 <= weights[3667];
				12'd3667	: data2 <= weights[3668];
				12'd3668	: data2 <= weights[3669];
				12'd3669	: data2 <= weights[3670];
				12'd3670	: data2 <= weights[3671];
				12'd3671	: data2 <= weights[3672];
				12'd3672	: data2 <= weights[3673];
				12'd3673	: data2 <= weights[3674];
				12'd3674	: data2 <= weights[3675];
				12'd3675	: data2 <= weights[3676];
				12'd3676	: data2 <= weights[3677];
				12'd3677	: data2 <= weights[3678];
				12'd3678	: data2 <= weights[3679];
				12'd3679	: data2 <= weights[3680];
				12'd3680	: data2 <= weights[3681];
				12'd3681	: data2 <= weights[3682];
				12'd3682	: data2 <= weights[3683];
				12'd3683	: data2 <= weights[3684];
				12'd3684	: data2 <= weights[3685];
				12'd3685	: data2 <= weights[3686];
				12'd3686	: data2 <= weights[3687];
				12'd3687	: data2 <= weights[3688];
				12'd3688	: data2 <= weights[3689];
				12'd3689	: data2 <= weights[3690];
				12'd3690	: data2 <= weights[3691];
				12'd3691	: data2 <= weights[3692];
				12'd3692	: data2 <= weights[3693];
				12'd3693	: data2 <= weights[3694];
				12'd3694	: data2 <= weights[3695];
				12'd3695	: data2 <= weights[3696];
				12'd3696	: data2 <= weights[3697];
				12'd3697	: data2 <= weights[3698];
				12'd3698	: data2 <= weights[3699];
				12'd3699	: data2 <= weights[3700];
				12'd3700	: data2 <= weights[3701];
				12'd3701	: data2 <= weights[3702];
				12'd3702	: data2 <= weights[3703];
				12'd3703	: data2 <= weights[3704];
				12'd3704	: data2 <= weights[3705];
				12'd3705	: data2 <= weights[3706];
				12'd3706	: data2 <= weights[3707];
				12'd3707	: data2 <= weights[3708];
				12'd3708	: data2 <= weights[3709];
				12'd3709	: data2 <= weights[3710];
				12'd3710	: data2 <= weights[3711];
				12'd3711	: data2 <= weights[3712];
				12'd3712	: data2 <= weights[3713];
				12'd3713	: data2 <= weights[3714];
				12'd3714	: data2 <= weights[3715];
				12'd3715	: data2 <= weights[3716];
				12'd3716	: data2 <= weights[3717];
				12'd3717	: data2 <= weights[3718];
				12'd3718	: data2 <= weights[3719];
				12'd3719	: data2 <= weights[3720];
				12'd3720	: data2 <= weights[3721];
				12'd3721	: data2 <= weights[3722];
				12'd3722	: data2 <= weights[3723];
				12'd3723	: data2 <= weights[3724];
				12'd3724	: data2 <= weights[3725];
				12'd3725	: data2 <= weights[3726];
				12'd3726	: data2 <= weights[3727];
				12'd3727	: data2 <= weights[3728];
				12'd3728	: data2 <= weights[3729];
				12'd3729	: data2 <= weights[3730];
				12'd3730	: data2 <= weights[3731];
				12'd3731	: data2 <= weights[3732];
				12'd3732	: data2 <= weights[3733];
				12'd3733	: data2 <= weights[3734];
				12'd3734	: data2 <= weights[3735];
				12'd3735	: data2 <= weights[3736];
				12'd3736	: data2 <= weights[3737];
				12'd3737	: data2 <= weights[3738];
				12'd3738	: data2 <= weights[3739];
				12'd3739	: data2 <= weights[3740];
				12'd3740	: data2 <= weights[3741];
				12'd3741	: data2 <= weights[3742];
				12'd3742	: data2 <= weights[3743];
				12'd3743	: data2 <= weights[3744];
				12'd3744	: data2 <= weights[3745];
				12'd3745	: data2 <= weights[3746];
				12'd3746	: data2 <= weights[3747];
				12'd3747	: data2 <= weights[3748];
				12'd3748	: data2 <= weights[3749];
				12'd3749	: data2 <= weights[3750];
				12'd3750	: data2 <= weights[3751];
				12'd3751	: data2 <= weights[3752];
				12'd3752	: data2 <= weights[3753];
				12'd3753	: data2 <= weights[3754];
				12'd3754	: data2 <= weights[3755];
				12'd3755	: data2 <= weights[3756];
				12'd3756	: data2 <= weights[3757];
				12'd3757	: data2 <= weights[3758];
				12'd3758	: data2 <= weights[3759];
				12'd3759	: data2 <= weights[3760];
				12'd3760	: data2 <= weights[3761];
				12'd3761	: data2 <= weights[3762];
				12'd3762	: data2 <= weights[3763];
				12'd3763	: data2 <= weights[3764];
				12'd3764	: data2 <= weights[3765];
				12'd3765	: data2 <= weights[3766];
				12'd3766	: data2 <= weights[3767];
				12'd3767	: data2 <= weights[3768];
				12'd3768	: data2 <= weights[3769];
				12'd3769	: data2 <= weights[3770];
				12'd3770	: data2 <= weights[3771];
				12'd3771	: data2 <= weights[3772];
				12'd3772	: data2 <= weights[3773];
				12'd3773	: data2 <= weights[3774];
				12'd3774	: data2 <= weights[3775];
				12'd3775	: data2 <= weights[3776];
				12'd3776	: data2 <= weights[3777];
				12'd3777	: data2 <= weights[3778];
				12'd3778	: data2 <= weights[3779];
				12'd3779	: data2 <= weights[3780];
				12'd3780	: data2 <= weights[3781];
				12'd3781	: data2 <= weights[3782];
				12'd3782	: data2 <= weights[3783];
				12'd3783	: data2 <= weights[3784];
				12'd3784	: data2 <= weights[3785];
				12'd3785	: data2 <= weights[3786];
				12'd3786	: data2 <= weights[3787];
				12'd3787	: data2 <= weights[3788];
				12'd3788	: data2 <= weights[3789];
				12'd3789	: data2 <= weights[3790];
				12'd3790	: data2 <= weights[3791];
				12'd3791	: data2 <= weights[3792];
				12'd3792	: data2 <= weights[3793];
				12'd3793	: data2 <= weights[3794];
				12'd3794	: data2 <= weights[3795];
				12'd3795	: data2 <= weights[3796];
				12'd3796	: data2 <= weights[3797];
				12'd3797	: data2 <= weights[3798];
				12'd3798	: data2 <= weights[3799];
				12'd3799	: data2 <= weights[3800];
				12'd3800	: data2 <= weights[3801];
				12'd3801	: data2 <= weights[3802];
				12'd3802	: data2 <= weights[3803];
				12'd3803	: data2 <= weights[3804];
				12'd3804	: data2 <= weights[3805];
				12'd3805	: data2 <= weights[3806];
				12'd3806	: data2 <= weights[3807];
				12'd3807	: data2 <= weights[3808];
				12'd3808	: data2 <= weights[3809];
				12'd3809	: data2 <= weights[3810];
				12'd3810	: data2 <= weights[3811];
				12'd3811	: data2 <= weights[3812];
				12'd3812	: data2 <= weights[3813];
				12'd3813	: data2 <= weights[3814];
				12'd3814	: data2 <= weights[3815];
				12'd3815	: data2 <= weights[3816];
				12'd3816	: data2 <= weights[3817];
				12'd3817	: data2 <= weights[3818];
				12'd3818	: data2 <= weights[3819];
				12'd3819	: data2 <= weights[3820];
				12'd3820	: data2 <= weights[3821];
				12'd3821	: data2 <= weights[3822];
				12'd3822	: data2 <= weights[3823];
				12'd3823	: data2 <= weights[3824];
				12'd3824	: data2 <= weights[3825];
				12'd3825	: data2 <= weights[3826];
				12'd3826	: data2 <= weights[3827];
				12'd3827	: data2 <= weights[3828];
				12'd3828	: data2 <= weights[3829];
				12'd3829	: data2 <= weights[3830];
				12'd3830	: data2 <= weights[3831];
				12'd3831	: data2 <= weights[3832];
				12'd3832	: data2 <= weights[3833];
				12'd3833	: data2 <= weights[3834];
				12'd3834	: data2 <= weights[3835];
				12'd3835	: data2 <= weights[3836];
				12'd3836	: data2 <= weights[3837];
				12'd3837	: data2 <= weights[3838];
				12'd3838	: data2 <= weights[3839];
				12'd3839	: data2 <= weights[3840];
				12'd3840	: data2 <= weights[3841];
				12'd3841	: data2 <= weights[3842];
				12'd3842	: data2 <= weights[3843];
				12'd3843	: data2 <= weights[3844];
				12'd3844	: data2 <= weights[3845];
				12'd3845	: data2 <= weights[3846];
				12'd3846	: data2 <= weights[3847];
				12'd3847	: data2 <= weights[3848];
				12'd3848	: data2 <= weights[3849];
				12'd3849	: data2 <= weights[3850];
				12'd3850	: data2 <= weights[3851];
				12'd3851	: data2 <= weights[3852];
				12'd3852	: data2 <= weights[3853];
				12'd3853	: data2 <= weights[3854];
				12'd3854	: data2 <= weights[3855];
				12'd3855	: data2 <= weights[3856];
				12'd3856	: data2 <= weights[3857];
				12'd3857	: data2 <= weights[3858];
				12'd3858	: data2 <= weights[3859];
				12'd3859	: data2 <= weights[3860];
				12'd3860	: data2 <= weights[3861];
				12'd3861	: data2 <= weights[3862];
				12'd3862	: data2 <= weights[3863];
				12'd3863	: data2 <= weights[3864];
				12'd3864	: data2 <= weights[3865];
				12'd3865	: data2 <= weights[3866];
				12'd3866	: data2 <= weights[3867];
				12'd3867	: data2 <= weights[3868];
				12'd3868	: data2 <= weights[3869];
				12'd3869	: data2 <= weights[3870];
				12'd3870	: data2 <= weights[3871];
				12'd3871	: data2 <= weights[3872];
				12'd3872	: data2 <= weights[3873];
				12'd3873	: data2 <= weights[3874];
				12'd3874	: data2 <= weights[3875];
				12'd3875	: data2 <= weights[3876];
				12'd3876	: data2 <= weights[3877];
				12'd3877	: data2 <= weights[3878];
				12'd3878	: data2 <= weights[3879];
				12'd3879	: data2 <= weights[3880];
				12'd3880	: data2 <= weights[3881];
				12'd3881	: data2 <= weights[3882];
				12'd3882	: data2 <= weights[3883];
				12'd3883	: data2 <= weights[3884];
				12'd3884	: data2 <= weights[3885];
				12'd3885	: data2 <= weights[3886];
				12'd3886	: data2 <= weights[3887];
				12'd3887	: data2 <= weights[3888];
				12'd3888	: data2 <= weights[3889];
				12'd3889	: data2 <= weights[3890];
				12'd3890	: data2 <= weights[3891];
				12'd3891	: data2 <= weights[3892];
				12'd3892	: data2 <= weights[3893];
				12'd3893	: data2 <= weights[3894];
				12'd3894	: data2 <= weights[3895];
				12'd3895	: data2 <= weights[3896];
				12'd3896	: data2 <= weights[3897];
				12'd3897	: data2 <= weights[3898];
				12'd3898	: data2 <= weights[3899];
				12'd3899	: data2 <= weights[3900];
				12'd3900	: data2 <= weights[3901];
				12'd3901	: data2 <= weights[3902];
				12'd3902	: data2 <= weights[3903];
				12'd3903	: data2 <= weights[3904];
				12'd3904	: data2 <= weights[3905];
				12'd3905	: data2 <= weights[3906];
				12'd3906	: data2 <= weights[3907];
				12'd3907	: data2 <= weights[3908];
				12'd3908	: data2 <= weights[3909];
				12'd3909	: data2 <= weights[3910];
				12'd3910	: data2 <= weights[3911];
				12'd3911	: data2 <= weights[3912];
				12'd3912	: data2 <= weights[3913];
				12'd3913	: data2 <= weights[3914];
				12'd3914	: data2 <= weights[3915];
				12'd3915	: data2 <= weights[3916];
				12'd3916	: data2 <= weights[3917];
				12'd3917	: data2 <= weights[3918];
				12'd3918	: data2 <= weights[3919];
				12'd3919	: data2 <= weights[3920];
				12'd3920	: data2 <= weights[3921];
				12'd3921	: data2 <= weights[3922];
				12'd3922	: data2 <= weights[3923];
				12'd3923	: data2 <= weights[3924];
				12'd3924	: data2 <= weights[3925];
				12'd3925	: data2 <= weights[3926];
				12'd3926	: data2 <= weights[3927];
				12'd3927	: data2 <= weights[3928];
				12'd3928	: data2 <= weights[3929];
				12'd3929	: data2 <= weights[3930];
				12'd3930	: data2 <= weights[3931];
				12'd3931	: data2 <= weights[3932];
				12'd3932	: data2 <= weights[3933];
				12'd3933	: data2 <= weights[3934];
				12'd3934	: data2 <= weights[3935];
				12'd3935	: data2 <= weights[3936];
				12'd3936	: data2 <= weights[3937];
				12'd3937	: data2 <= weights[3938];
				12'd3938	: data2 <= weights[3939];
				12'd3939	: data2 <= weights[3940];
				12'd3940	: data2 <= weights[3941];
				12'd3941	: data2 <= weights[3942];
				12'd3942	: data2 <= weights[3943];
				12'd3943	: data2 <= weights[3944];
				12'd3944	: data2 <= weights[3945];
				12'd3945	: data2 <= weights[3946];
				12'd3946	: data2 <= weights[3947];
				12'd3947	: data2 <= weights[3948];
				12'd3948	: data2 <= weights[3949];
				12'd3949	: data2 <= weights[3950];
				12'd3950	: data2 <= weights[3951];
				12'd3951	: data2 <= weights[3952];
				12'd3952	: data2 <= weights[3953];
				12'd3953	: data2 <= weights[3954];
				12'd3954	: data2 <= weights[3955];
				12'd3955	: data2 <= weights[3956];
				12'd3956	: data2 <= weights[3957];
				12'd3957	: data2 <= weights[3958];
				12'd3958	: data2 <= weights[3959];
				12'd3959	: data2 <= weights[3960];
				12'd3960	: data2 <= weights[3961];
				12'd3961	: data2 <= weights[3962];
				12'd3962	: data2 <= weights[3963];
				12'd3963	: data2 <= weights[3964];
				12'd3964	: data2 <= weights[3965];
				12'd3965	: data2 <= weights[3966];
				12'd3966	: data2 <= weights[3967];
				12'd3967	: data2 <= weights[3968];
				12'd3968	: data2 <= weights[3969];
				12'd3969	: data2 <= weights[3970];
				12'd3970	: data2 <= weights[3971];
				12'd3971	: data2 <= weights[3972];
				12'd3972	: data2 <= weights[3973];
				12'd3973	: data2 <= weights[3974];
				12'd3974	: data2 <= weights[3975];
				12'd3975	: data2 <= weights[3976];
				12'd3976	: data2 <= weights[3977];
				12'd3977	: data2 <= weights[3978];
				12'd3978	: data2 <= weights[3979];
				12'd3979	: data2 <= weights[3980];
				12'd3980	: data2 <= weights[3981];
				12'd3981	: data2 <= weights[3982];
				12'd3982	: data2 <= weights[3983];
				12'd3983	: data2 <= weights[3984];
				12'd3984	: data2 <= weights[3985];
				12'd3985	: data2 <= weights[3986];
				12'd3986	: data2 <= weights[3987];
				12'd3987	: data2 <= weights[3988];
				12'd3988	: data2 <= weights[3989];
				12'd3989	: data2 <= weights[3990];
				12'd3990	: data2 <= weights[3991];
				12'd3991	: data2 <= weights[3992];
				12'd3992	: data2 <= weights[3993];
				12'd3993	: data2 <= weights[3994];
				12'd3994	: data2 <= weights[3995];
				12'd3995	: data2 <= weights[3996];
				12'd3996	: data2 <= weights[3997];
				12'd3997	: data2 <= weights[3998];
				12'd3998	: data2 <= weights[3999];
				12'd3999	: data2 <= weights[4000];
				12'd4000	: data2 <= weights[4001];
				12'd4001	: data2 <= weights[4002];
				12'd4002	: data2 <= weights[4003];
				12'd4003	: data2 <= weights[4004];
				12'd4004	: data2 <= weights[4005];
				12'd4005	: data2 <= weights[4006];
				12'd4006	: data2 <= weights[4007];
				12'd4007	: data2 <= weights[4008];
				12'd4008	: data2 <= weights[4009];
				12'd4009	: data2 <= weights[4010];
				12'd4010	: data2 <= weights[4011];
				12'd4011	: data2 <= weights[4012];
				12'd4012	: data2 <= weights[4013];
				12'd4013	: data2 <= weights[4014];
				12'd4014	: data2 <= weights[4015];
				12'd4015	: data2 <= weights[4016];
				12'd4016	: data2 <= weights[4017];
				12'd4017	: data2 <= weights[4018];
				12'd4018	: data2 <= weights[4019];
				12'd4019	: data2 <= weights[4020];
				12'd4020	: data2 <= weights[4021];
				12'd4021	: data2 <= weights[4022];
				12'd4022	: data2 <= weights[4023];
				12'd4023	: data2 <= weights[4024];
				12'd4024	: data2 <= weights[4025];
				12'd4025	: data2 <= weights[4026];
				12'd4026	: data2 <= weights[4027];
				12'd4027	: data2 <= weights[4028];
				12'd4028	: data2 <= weights[4029];
				12'd4029	: data2 <= weights[4030];
				12'd4030	: data2 <= weights[4031];
				12'd4031	: data2 <= weights[4032];
				12'd4032	: data2 <= weights[4033];
				12'd4033	: data2 <= weights[4034];
				12'd4034	: data2 <= weights[4035];
				12'd4035	: data2 <= weights[4036];
				12'd4036	: data2 <= weights[4037];
				12'd4037	: data2 <= weights[4038];
				12'd4038	: data2 <= weights[4039];
				12'd4039	: data2 <= weights[4040];
				12'd4040	: data2 <= weights[4041];
				12'd4041	: data2 <= weights[4042];
				12'd4042	: data2 <= weights[4043];
				12'd4043	: data2 <= weights[4044];
				12'd4044	: data2 <= weights[4045];
				12'd4045	: data2 <= weights[4046];
				12'd4046	: data2 <= weights[4047];
				12'd4047	: data2 <= weights[4048];
				12'd4048	: data2 <= weights[4049];
				12'd4049	: data2 <= weights[4050];
				default		: data2 <= 16'd0;
			endcase
		end else begin
			data2 <= data2;
		end
	end

endmodule