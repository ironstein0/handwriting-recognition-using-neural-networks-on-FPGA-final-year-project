`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   09:00:54 02/26/2016
// Design Name:   sigmoid
// Module Name:   /home/kishore/Desktop/verilog_files/final_sigmoid_try/sigmoid_tb.v
// Project Name:  final_sigmoid_try
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: sigmoid
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module sigmoid_tb;

	// Inputs
	reg clk;
	reg reset;
	reg [17:0] x1;
	//real itr=-5.0;
	//real tmp;

	// Outputs
	wire [47:0] fixed_op;
//	wire [2:0] test;
	// Instantiate the Unit Under Test (UUT)
	sigmoid uut (
		.clk(clk), 
		.reset(reset),
		.x1(x1), 
		.fixed_op(fixed_op)
//		.test(test)
	);

	always begin
		#1 clk = ~ clk;
	end

	initial begin
		// Initialize Inputs
		clk = 0;
		//-11.0
		#61
		x1=18'b1_1011_0000000000000;
		
		//-10.6
		#60
		x1=18'b1_1010_1001100110011;

		//-10.2
		#60
		x1=18'b1_1010_0011001100110;

		//-9.8
		#60
		x1=18'b1_1001_1100110011010;

		//-9.4
		#60
		x1=18'b1_1001_0110011001101;

		//-9.0
		#60
		x1=18'b1_1001_0000000000000;

		//-8.6
		#60
		x1=18'b1_1000_1001100110011;

		//-8.2
		#60
		x1=18'b1_1000_0011001100110;

		//-7.8
		#60
		x1=18'b1_0111_1100110011010;

		//-7.4
		#60
		x1=18'b1_0111_0110011001101;

		//-7.0
		#60
		x1=18'b1_0111_1000000000000;

		//-6.6
		#60
		x1=18'b1_0110_1001100110011;

		//-6.2
		#60
		x1=18'b1_0110_0011001100110;

		//-5.8
		#60
		x1=18'b1_0101_1100110011010;

		//-5.4
		#60
		x1=18'b1_0101_0110011001101;

		//-5.0
		#60
		x1=18'b1_0101_0000000000000;

		//-4.6
		#60
		x1=18'b1_0100_1001100110011;

		//-4.2
		#60
		x1=18'b1_0100_0011001100110;

		//-3.8
		#60
		x1=18'b1_0011_1100110011010;

		//-3.4
		#60
		x1=18'b1_0011_0110011001101;

		//-3.0
		#60
		x1=18'b1_0011_0000000000000;

		//-2.6
		#60
		x1=18'b1_0010_1001100110011;

		//-2.2
		#60
		x1=18'b1_0010_0011001100110;

		//-1.8
		#60
		x1=18'b1_0001_1100110011010;

		//-1.4
		#60
		x1=18'b1_0001_0110011001101;

		//-1.0
		#60
		x1=18'b1_0001_0000000000000;

		//-0.6
		#60
		x1=18'b1_0000_1001100110011;

		//-0.2
		#60
		x1=18'b1_0000_0011001100110;

		//0.2
		#60
		x1=18'b0_0000_0011001100110;

		//0.6
		#60
		x1=18'b0_0000_1001100110011;

		//1.0
		#60
		x1=18'b0_0001_0000000000000;

		//1.4
		#60
		x1=18'b0_0001_0110011001101;

		//1.8
		#60
		x1=18'b0_0001_1100110011010;

		//2.2
		#60
		x1=18'b0_0010_0011001100110;

		//2.6
		#60
		x1=18'b0_0010_1001100110011;

		//3.0
		#60
		x1=18'b0_0011_0000000000000;

		//3.4
		#60
		x1=18'b0_0011_0110011001101;

		//3.8
		#60
		x1=18'b0_0011_1100110011010;

		//4.2
		#60
		x1=18'b0_0100_0011001100110;

		//4.6
		#60
		x1=18'b0_0100_1001100110011;

		//5.0
		#60
		x1=18'b0_0101_0000000000000;

		//5.4
		#60
		x1=18'b0_0101_0110011001101;

		//5.8
		#60
		x1=18'b0_0101_1100110011010;

		//6.2
		#60
		x1=18'b0_0110_0011001100110;

		//6.6
		#60
		x1=18'b0_0110_1001100110011;

		//7.0
		#60
		x1=18'b0_0111_0000000000000;

		//7.4
		#60
		x1=18'b0_0111_0110011001101;

		//7.8
		#60
		x1=18'b0_0111_1100110011010;

		//8.2
		#60
		x1=18'b0_1000_0011001100110;

		//8.6
		#60
		x1=18'b0_1000_1001100110011;

		//9.0
		#60
		x1=18'b0_1001_0000000000000;

		//9.4
		#60
		x1=18'b0_1001_0110011001101;

		//9.8
		#60
		x1=18'b0_1001_1100110011010;

		//10.2
		#60
		x1=18'b0_1010_0011001100110;

		//10.6
		#60
		x1=18'b0_1010_1001100110011;

		//11.0
		#60
		x1=18'b0_1011_0000000000000;
		
		#11 reset = 1;
		#10 reset = 0;

	end
/********this code works,DO NOT CHANGE********/		
		//$dumpfile("/home/kishore/Desktop/sigmoid_plot.vcd");
		//$dumpvars(1,x,fixed_op);//plot only changes in x and fixed_op
		//$dumpoff;
		// Wait 100 ns for global reset to finish
		
        
		// Add stimulus here
		//fixed_op takes at least two clock cycles
//		#40
//		//x=18'b00100_1111111110111;    binary
//		 //$dumpon;
//		 x=18'h09ff7;               // or hex format of +4.999
//		 //$dumpoff;
//		#40
//		//x=18'b00110_0001100110011;//+6.1
//		//$dumpon;
//		x=18'hc333;
//		//$dumpoff;
//		#40
//		//x=18'b00010_1100110011001;//+2.8
//		//$dumpon ;
//		x=18'h5999;
//		//$dumpoff;
//		#40
//		//x=18'b00000_1110000000000;//+0.875
//		//$dumpon;
//		x=18'h1c00;
//		end
//		//$dumpoff;
	initial begin
		$monitor("x: %h  ,fixed_op:%d",x1,fixed_op);
	end
	
	
//	always begin
//	#20 clk=~clk;
//	end
      
endmodule

