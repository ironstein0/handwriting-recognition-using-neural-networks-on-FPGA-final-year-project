module main;
initial
	begin
		$display("learning verilog is very easy");
		$finish;
	end
endmodule