`timescale 1ns / 1ps
`include "seven_segment_display_controller.v"
`include "binary_to_12bit_bcd_converter.v"
module stimulus(
    );


endmodule
